
module rca_N32 ( A, B, S, Co );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  output Co;
  wire   \CTMP[9] , \CTMP[8] , \CTMP[7] , \CTMP[6] , \CTMP[5] , \CTMP[4] ,
         \CTMP[3] , \CTMP[31] , \CTMP[30] , \CTMP[2] , \CTMP[29] , \CTMP[28] ,
         \CTMP[27] , \CTMP[26] , \CTMP[25] , \CTMP[24] , \CTMP[23] ,
         \CTMP[22] , \CTMP[21] , \CTMP[20] , \CTMP[1] , \CTMP[19] , \CTMP[18] ,
         \CTMP[17] , \CTMP[16] , \CTMP[15] , \CTMP[14] , \CTMP[13] ,
         \CTMP[12] , \CTMP[11] , \CTMP[10] ;

  HA_1 HA_0 ( .A(A[0]), .B(B[0]), .S(S[0]), .Co(\CTMP[1] ) );
  FA_159 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(\CTMP[1] ), .S(S[1]), .Co(\CTMP[2] )
         );
  FA_158 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(\CTMP[2] ), .S(S[2]), .Co(\CTMP[3] )
         );
  FA_157 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(\CTMP[3] ), .S(S[3]), .Co(\CTMP[4] )
         );
  FA_156 FA_i_5 ( .A(A[4]), .B(B[4]), .Ci(\CTMP[4] ), .S(S[4]), .Co(\CTMP[5] )
         );
  FA_155 FA_i_6 ( .A(A[5]), .B(B[5]), .Ci(\CTMP[5] ), .S(S[5]), .Co(\CTMP[6] )
         );
  FA_154 FA_i_7 ( .A(A[6]), .B(B[6]), .Ci(\CTMP[6] ), .S(S[6]), .Co(\CTMP[7] )
         );
  FA_153 FA_i_8 ( .A(A[7]), .B(B[7]), .Ci(\CTMP[7] ), .S(S[7]), .Co(\CTMP[8] )
         );
  FA_152 FA_i_9 ( .A(A[8]), .B(B[8]), .Ci(\CTMP[8] ), .S(S[8]), .Co(\CTMP[9] )
         );
  FA_151 FA_i_10 ( .A(A[9]), .B(B[9]), .Ci(\CTMP[9] ), .S(S[9]), .Co(
        \CTMP[10] ) );
  FA_150 FA_i_11 ( .A(A[10]), .B(B[10]), .Ci(\CTMP[10] ), .S(S[10]), .Co(
        \CTMP[11] ) );
  FA_149 FA_i_12 ( .A(A[11]), .B(B[11]), .Ci(\CTMP[11] ), .S(S[11]), .Co(
        \CTMP[12] ) );
  FA_148 FA_i_13 ( .A(A[12]), .B(B[12]), .Ci(\CTMP[12] ), .S(S[12]), .Co(
        \CTMP[13] ) );
  FA_147 FA_i_14 ( .A(A[13]), .B(B[13]), .Ci(\CTMP[13] ), .S(S[13]), .Co(
        \CTMP[14] ) );
  FA_146 FA_i_15 ( .A(A[14]), .B(B[14]), .Ci(\CTMP[14] ), .S(S[14]), .Co(
        \CTMP[15] ) );
  FA_145 FA_i_16 ( .A(A[15]), .B(B[15]), .Ci(\CTMP[15] ), .S(S[15]), .Co(
        \CTMP[16] ) );
  FA_144 FA_i_17 ( .A(A[16]), .B(B[16]), .Ci(\CTMP[16] ), .S(S[16]), .Co(
        \CTMP[17] ) );
  FA_143 FA_i_18 ( .A(A[17]), .B(B[17]), .Ci(\CTMP[17] ), .S(S[17]), .Co(
        \CTMP[18] ) );
  FA_142 FA_i_19 ( .A(A[18]), .B(B[18]), .Ci(\CTMP[18] ), .S(S[18]), .Co(
        \CTMP[19] ) );
  FA_141 FA_i_20 ( .A(A[19]), .B(B[19]), .Ci(\CTMP[19] ), .S(S[19]), .Co(
        \CTMP[20] ) );
  FA_140 FA_i_21 ( .A(A[20]), .B(B[20]), .Ci(\CTMP[20] ), .S(S[20]), .Co(
        \CTMP[21] ) );
  FA_139 FA_i_22 ( .A(A[21]), .B(B[21]), .Ci(\CTMP[21] ), .S(S[21]), .Co(
        \CTMP[22] ) );
  FA_138 FA_i_23 ( .A(A[22]), .B(B[22]), .Ci(\CTMP[22] ), .S(S[22]), .Co(
        \CTMP[23] ) );
  FA_137 FA_i_24 ( .A(A[23]), .B(B[23]), .Ci(\CTMP[23] ), .S(S[23]), .Co(
        \CTMP[24] ) );
  FA_136 FA_i_25 ( .A(A[24]), .B(B[24]), .Ci(\CTMP[24] ), .S(S[24]), .Co(
        \CTMP[25] ) );
  FA_135 FA_i_26 ( .A(A[25]), .B(B[25]), .Ci(\CTMP[25] ), .S(S[25]), .Co(
        \CTMP[26] ) );
  FA_134 FA_i_27 ( .A(A[26]), .B(B[26]), .Ci(\CTMP[26] ), .S(S[26]), .Co(
        \CTMP[27] ) );
  FA_133 FA_i_28 ( .A(A[27]), .B(B[27]), .Ci(\CTMP[27] ), .S(S[27]), .Co(
        \CTMP[28] ) );
  FA_132 FA_i_29 ( .A(A[28]), .B(B[28]), .Ci(\CTMP[28] ), .S(S[28]), .Co(
        \CTMP[29] ) );
  FA_131 FA_i_30 ( .A(A[29]), .B(B[29]), .Ci(\CTMP[29] ), .S(S[29]), .Co(
        \CTMP[30] ) );
  FA_130 FA_i_31 ( .A(A[30]), .B(B[30]), .Ci(\CTMP[30] ), .S(S[30]), .Co(
        \CTMP[31] ) );
  FA_129 FA_i_32 ( .A(A[31]), .B(B[31]), .Ci(\CTMP[31] ), .S(S[31]), .Co(Co)
         );
endmodule


module mux5to1_N32 ( A, B, C, D, E, Y, SEL );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  output [31:0] Y;
  input [2:0] SEL;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314;

  BUF_X1 U1 ( .A(n9), .Z(n302) );
  BUF_X1 U2 ( .A(n8), .Z(n304) );
  BUF_X1 U3 ( .A(n8), .Z(n303) );
  BUF_X1 U4 ( .A(n9), .Z(n301) );
  BUF_X1 U5 ( .A(n9), .Z(n300) );
  BUF_X1 U6 ( .A(n6), .Z(n310) );
  BUF_X1 U7 ( .A(n6), .Z(n309) );
  BUF_X1 U8 ( .A(n7), .Z(n307) );
  BUF_X1 U9 ( .A(n7), .Z(n306) );
  BUF_X1 U10 ( .A(n5), .Z(n313) );
  BUF_X1 U11 ( .A(n5), .Z(n312) );
  BUF_X1 U12 ( .A(n8), .Z(n305) );
  BUF_X1 U13 ( .A(n6), .Z(n311) );
  BUF_X1 U14 ( .A(n7), .Z(n308) );
  BUF_X1 U15 ( .A(n5), .Z(n314) );
  NOR3_X1 U16 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n72), .ZN(n6) );
  NOR3_X1 U17 ( .A1(n72), .A2(SEL[2]), .A3(n73), .ZN(n7) );
  NOR3_X1 U18 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n73), .ZN(n8) );
  NOR2_X1 U19 ( .A1(n74), .A2(n302), .ZN(n5) );
  AOI21_X1 U20 ( .B1(n72), .B2(n73), .A(SEL[2]), .ZN(n74) );
  INV_X1 U21 ( .A(SEL[0]), .ZN(n73) );
  INV_X1 U22 ( .A(SEL[1]), .ZN(n72) );
  AND3_X1 U23 ( .A1(n73), .A2(n72), .A3(SEL[2]), .ZN(n9) );
  NAND2_X1 U24 ( .A1(n22), .A2(n23), .ZN(Y[31]) );
  AOI22_X1 U25 ( .A1(B[31]), .A2(n305), .B1(E[31]), .B2(n300), .ZN(n22) );
  AOI222_X1 U26 ( .A1(A[31]), .A2(n314), .B1(C[31]), .B2(n311), .C1(D[31]), 
        .C2(n308), .ZN(n23) );
  NAND2_X1 U27 ( .A1(n3), .A2(n4), .ZN(Y[9]) );
  AOI22_X1 U28 ( .A1(B[9]), .A2(n305), .B1(E[9]), .B2(n301), .ZN(n3) );
  AOI222_X1 U29 ( .A1(A[9]), .A2(n314), .B1(C[9]), .B2(n311), .C1(D[9]), .C2(
        n308), .ZN(n4) );
  NAND2_X1 U30 ( .A1(n10), .A2(n11), .ZN(Y[8]) );
  AOI22_X1 U31 ( .A1(B[8]), .A2(n305), .B1(E[8]), .B2(n300), .ZN(n10) );
  AOI222_X1 U32 ( .A1(A[8]), .A2(n314), .B1(C[8]), .B2(n311), .C1(D[8]), .C2(
        n308), .ZN(n11) );
  NAND2_X1 U33 ( .A1(n12), .A2(n13), .ZN(Y[7]) );
  AOI22_X1 U34 ( .A1(B[7]), .A2(n305), .B1(E[7]), .B2(n300), .ZN(n12) );
  AOI222_X1 U35 ( .A1(A[7]), .A2(n314), .B1(C[7]), .B2(n311), .C1(D[7]), .C2(
        n308), .ZN(n13) );
  NAND2_X1 U36 ( .A1(n14), .A2(n15), .ZN(Y[6]) );
  AOI22_X1 U37 ( .A1(B[6]), .A2(n305), .B1(E[6]), .B2(n300), .ZN(n14) );
  AOI222_X1 U38 ( .A1(A[6]), .A2(n314), .B1(C[6]), .B2(n311), .C1(D[6]), .C2(
        n308), .ZN(n15) );
  NAND2_X1 U39 ( .A1(n16), .A2(n17), .ZN(Y[5]) );
  AOI22_X1 U40 ( .A1(B[5]), .A2(n305), .B1(E[5]), .B2(n300), .ZN(n16) );
  AOI222_X1 U41 ( .A1(A[5]), .A2(n314), .B1(C[5]), .B2(n311), .C1(D[5]), .C2(
        n308), .ZN(n17) );
  NAND2_X1 U42 ( .A1(n18), .A2(n19), .ZN(Y[4]) );
  AOI22_X1 U43 ( .A1(B[4]), .A2(n305), .B1(E[4]), .B2(n300), .ZN(n18) );
  AOI222_X1 U44 ( .A1(A[4]), .A2(n314), .B1(C[4]), .B2(n311), .C1(D[4]), .C2(
        n308), .ZN(n19) );
  NAND2_X1 U45 ( .A1(n20), .A2(n21), .ZN(Y[3]) );
  AOI22_X1 U46 ( .A1(B[3]), .A2(n305), .B1(E[3]), .B2(n300), .ZN(n20) );
  AOI222_X1 U47 ( .A1(A[3]), .A2(n314), .B1(C[3]), .B2(n311), .C1(D[3]), .C2(
        n308), .ZN(n21) );
  NAND2_X1 U48 ( .A1(n24), .A2(n25), .ZN(Y[30]) );
  AOI22_X1 U49 ( .A1(B[30]), .A2(n304), .B1(E[30]), .B2(n300), .ZN(n24) );
  AOI222_X1 U50 ( .A1(A[30]), .A2(n313), .B1(C[30]), .B2(n310), .C1(D[30]), 
        .C2(n307), .ZN(n25) );
  NAND2_X1 U51 ( .A1(n28), .A2(n29), .ZN(Y[29]) );
  AOI22_X1 U52 ( .A1(B[29]), .A2(n304), .B1(E[29]), .B2(n300), .ZN(n28) );
  AOI222_X1 U53 ( .A1(A[29]), .A2(n313), .B1(C[29]), .B2(n310), .C1(D[29]), 
        .C2(n307), .ZN(n29) );
  NAND2_X1 U54 ( .A1(n30), .A2(n31), .ZN(Y[28]) );
  AOI22_X1 U55 ( .A1(B[28]), .A2(n304), .B1(E[28]), .B2(n300), .ZN(n30) );
  AOI222_X1 U56 ( .A1(A[28]), .A2(n313), .B1(C[28]), .B2(n310), .C1(D[28]), 
        .C2(n307), .ZN(n31) );
  NAND2_X1 U57 ( .A1(n32), .A2(n33), .ZN(Y[27]) );
  AOI22_X1 U58 ( .A1(B[27]), .A2(n304), .B1(E[27]), .B2(n301), .ZN(n32) );
  AOI222_X1 U59 ( .A1(A[27]), .A2(n313), .B1(C[27]), .B2(n310), .C1(D[27]), 
        .C2(n307), .ZN(n33) );
  NAND2_X1 U60 ( .A1(n34), .A2(n35), .ZN(Y[26]) );
  AOI22_X1 U61 ( .A1(B[26]), .A2(n304), .B1(E[26]), .B2(n301), .ZN(n34) );
  AOI222_X1 U62 ( .A1(A[26]), .A2(n313), .B1(C[26]), .B2(n310), .C1(D[26]), 
        .C2(n307), .ZN(n35) );
  NAND2_X1 U63 ( .A1(n36), .A2(n37), .ZN(Y[25]) );
  AOI22_X1 U64 ( .A1(B[25]), .A2(n304), .B1(E[25]), .B2(n301), .ZN(n36) );
  AOI222_X1 U65 ( .A1(A[25]), .A2(n313), .B1(C[25]), .B2(n310), .C1(D[25]), 
        .C2(n307), .ZN(n37) );
  NAND2_X1 U66 ( .A1(n38), .A2(n39), .ZN(Y[24]) );
  AOI22_X1 U67 ( .A1(B[24]), .A2(n304), .B1(E[24]), .B2(n301), .ZN(n38) );
  AOI222_X1 U68 ( .A1(A[24]), .A2(n313), .B1(C[24]), .B2(n310), .C1(D[24]), 
        .C2(n307), .ZN(n39) );
  NAND2_X1 U69 ( .A1(n40), .A2(n41), .ZN(Y[23]) );
  AOI22_X1 U70 ( .A1(B[23]), .A2(n304), .B1(E[23]), .B2(n301), .ZN(n40) );
  AOI222_X1 U71 ( .A1(A[23]), .A2(n313), .B1(C[23]), .B2(n310), .C1(D[23]), 
        .C2(n307), .ZN(n41) );
  NAND2_X1 U72 ( .A1(n42), .A2(n43), .ZN(Y[22]) );
  AOI22_X1 U73 ( .A1(B[22]), .A2(n304), .B1(E[22]), .B2(n301), .ZN(n42) );
  AOI222_X1 U74 ( .A1(A[22]), .A2(n313), .B1(C[22]), .B2(n310), .C1(D[22]), 
        .C2(n307), .ZN(n43) );
  NAND2_X1 U75 ( .A1(n44), .A2(n45), .ZN(Y[21]) );
  AOI22_X1 U76 ( .A1(B[21]), .A2(n304), .B1(E[21]), .B2(n301), .ZN(n44) );
  AOI222_X1 U77 ( .A1(A[21]), .A2(n313), .B1(C[21]), .B2(n310), .C1(D[21]), 
        .C2(n307), .ZN(n45) );
  NAND2_X1 U78 ( .A1(n46), .A2(n47), .ZN(Y[20]) );
  AOI22_X1 U79 ( .A1(B[20]), .A2(n304), .B1(E[20]), .B2(n301), .ZN(n46) );
  AOI222_X1 U80 ( .A1(A[20]), .A2(n313), .B1(C[20]), .B2(n310), .C1(D[20]), 
        .C2(n307), .ZN(n47) );
  NAND2_X1 U81 ( .A1(n50), .A2(n51), .ZN(Y[19]) );
  AOI22_X1 U82 ( .A1(B[19]), .A2(n303), .B1(E[19]), .B2(n301), .ZN(n50) );
  AOI222_X1 U83 ( .A1(A[19]), .A2(n312), .B1(C[19]), .B2(n309), .C1(D[19]), 
        .C2(n306), .ZN(n51) );
  NAND2_X1 U84 ( .A1(n52), .A2(n53), .ZN(Y[18]) );
  AOI22_X1 U85 ( .A1(B[18]), .A2(n303), .B1(E[18]), .B2(n301), .ZN(n52) );
  AOI222_X1 U86 ( .A1(A[18]), .A2(n312), .B1(C[18]), .B2(n309), .C1(D[18]), 
        .C2(n306), .ZN(n53) );
  NAND2_X1 U87 ( .A1(n54), .A2(n55), .ZN(Y[17]) );
  AOI22_X1 U88 ( .A1(B[17]), .A2(n303), .B1(E[17]), .B2(n302), .ZN(n54) );
  AOI222_X1 U89 ( .A1(A[17]), .A2(n312), .B1(C[17]), .B2(n309), .C1(D[17]), 
        .C2(n306), .ZN(n55) );
  NAND2_X1 U90 ( .A1(n56), .A2(n57), .ZN(Y[16]) );
  AOI22_X1 U91 ( .A1(B[16]), .A2(n303), .B1(E[16]), .B2(n302), .ZN(n56) );
  AOI222_X1 U92 ( .A1(A[16]), .A2(n312), .B1(C[16]), .B2(n309), .C1(D[16]), 
        .C2(n306), .ZN(n57) );
  NAND2_X1 U93 ( .A1(n58), .A2(n59), .ZN(Y[15]) );
  AOI22_X1 U94 ( .A1(B[15]), .A2(n303), .B1(E[15]), .B2(n302), .ZN(n58) );
  AOI222_X1 U95 ( .A1(A[15]), .A2(n312), .B1(C[15]), .B2(n309), .C1(D[15]), 
        .C2(n306), .ZN(n59) );
  NAND2_X1 U96 ( .A1(n60), .A2(n61), .ZN(Y[14]) );
  AOI22_X1 U97 ( .A1(B[14]), .A2(n303), .B1(E[14]), .B2(n302), .ZN(n60) );
  AOI222_X1 U98 ( .A1(A[14]), .A2(n312), .B1(C[14]), .B2(n309), .C1(D[14]), 
        .C2(n306), .ZN(n61) );
  NAND2_X1 U99 ( .A1(n62), .A2(n63), .ZN(Y[13]) );
  AOI22_X1 U100 ( .A1(B[13]), .A2(n303), .B1(E[13]), .B2(n302), .ZN(n62) );
  AOI222_X1 U101 ( .A1(A[13]), .A2(n312), .B1(C[13]), .B2(n309), .C1(D[13]), 
        .C2(n306), .ZN(n63) );
  NAND2_X1 U102 ( .A1(n64), .A2(n65), .ZN(Y[12]) );
  AOI22_X1 U103 ( .A1(B[12]), .A2(n303), .B1(E[12]), .B2(n302), .ZN(n64) );
  AOI222_X1 U104 ( .A1(A[12]), .A2(n312), .B1(C[12]), .B2(n309), .C1(D[12]), 
        .C2(n306), .ZN(n65) );
  NAND2_X1 U105 ( .A1(n66), .A2(n67), .ZN(Y[11]) );
  AOI22_X1 U106 ( .A1(B[11]), .A2(n303), .B1(E[11]), .B2(n302), .ZN(n66) );
  AOI222_X1 U107 ( .A1(A[11]), .A2(n312), .B1(C[11]), .B2(n309), .C1(D[11]), 
        .C2(n306), .ZN(n67) );
  NAND2_X1 U108 ( .A1(n68), .A2(n69), .ZN(Y[10]) );
  AOI22_X1 U109 ( .A1(B[10]), .A2(n303), .B1(E[10]), .B2(n302), .ZN(n68) );
  AOI222_X1 U110 ( .A1(A[10]), .A2(n312), .B1(C[10]), .B2(n309), .C1(D[10]), 
        .C2(n306), .ZN(n69) );
  NAND2_X1 U111 ( .A1(n26), .A2(n27), .ZN(Y[2]) );
  AOI22_X1 U112 ( .A1(B[2]), .A2(n304), .B1(E[2]), .B2(n300), .ZN(n26) );
  AOI222_X1 U113 ( .A1(A[2]), .A2(n313), .B1(C[2]), .B2(n310), .C1(D[2]), .C2(
        n307), .ZN(n27) );
  NAND2_X1 U114 ( .A1(n48), .A2(n49), .ZN(Y[1]) );
  AOI22_X1 U115 ( .A1(B[1]), .A2(n303), .B1(E[1]), .B2(n301), .ZN(n48) );
  AOI222_X1 U116 ( .A1(A[1]), .A2(n312), .B1(C[1]), .B2(n309), .C1(D[1]), .C2(
        n306), .ZN(n49) );
  NAND2_X1 U117 ( .A1(n70), .A2(n71), .ZN(Y[0]) );
  AOI22_X1 U118 ( .A1(B[0]), .A2(n303), .B1(E[0]), .B2(n300), .ZN(n70) );
  AOI222_X1 U119 ( .A1(A[0]), .A2(n312), .B1(C[0]), .B2(n309), .C1(D[0]), .C2(
        n306), .ZN(n71) );
endmodule


module rca_N30 ( A, B, S, Co );
  input [29:0] A;
  input [29:0] B;
  output [29:0] S;
  output Co;
  wire   \CTMP[9] , \CTMP[8] , \CTMP[7] , \CTMP[6] , \CTMP[5] , \CTMP[4] ,
         \CTMP[3] , \CTMP[2] , \CTMP[29] , \CTMP[28] , \CTMP[27] , \CTMP[26] ,
         \CTMP[25] , \CTMP[24] , \CTMP[23] , \CTMP[22] , \CTMP[21] ,
         \CTMP[20] , \CTMP[1] , \CTMP[19] , \CTMP[18] , \CTMP[17] , \CTMP[16] ,
         \CTMP[15] , \CTMP[14] , \CTMP[13] , \CTMP[12] , \CTMP[11] ,
         \CTMP[10] ;

  HA_2 HA_0 ( .A(A[0]), .B(B[0]), .S(S[0]), .Co(\CTMP[1] ) );
  FA_188 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(\CTMP[1] ), .S(S[1]), .Co(\CTMP[2] )
         );
  FA_187 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(\CTMP[2] ), .S(S[2]), .Co(\CTMP[3] )
         );
  FA_186 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(\CTMP[3] ), .S(S[3]), .Co(\CTMP[4] )
         );
  FA_185 FA_i_5 ( .A(A[4]), .B(B[4]), .Ci(\CTMP[4] ), .S(S[4]), .Co(\CTMP[5] )
         );
  FA_184 FA_i_6 ( .A(A[5]), .B(B[5]), .Ci(\CTMP[5] ), .S(S[5]), .Co(\CTMP[6] )
         );
  FA_183 FA_i_7 ( .A(A[6]), .B(B[6]), .Ci(\CTMP[6] ), .S(S[6]), .Co(\CTMP[7] )
         );
  FA_182 FA_i_8 ( .A(A[7]), .B(B[7]), .Ci(\CTMP[7] ), .S(S[7]), .Co(\CTMP[8] )
         );
  FA_181 FA_i_9 ( .A(A[8]), .B(B[8]), .Ci(\CTMP[8] ), .S(S[8]), .Co(\CTMP[9] )
         );
  FA_180 FA_i_10 ( .A(A[9]), .B(B[9]), .Ci(\CTMP[9] ), .S(S[9]), .Co(
        \CTMP[10] ) );
  FA_179 FA_i_11 ( .A(A[10]), .B(B[10]), .Ci(\CTMP[10] ), .S(S[10]), .Co(
        \CTMP[11] ) );
  FA_178 FA_i_12 ( .A(A[11]), .B(B[11]), .Ci(\CTMP[11] ), .S(S[11]), .Co(
        \CTMP[12] ) );
  FA_177 FA_i_13 ( .A(A[12]), .B(B[12]), .Ci(\CTMP[12] ), .S(S[12]), .Co(
        \CTMP[13] ) );
  FA_176 FA_i_14 ( .A(A[13]), .B(B[13]), .Ci(\CTMP[13] ), .S(S[13]), .Co(
        \CTMP[14] ) );
  FA_175 FA_i_15 ( .A(A[14]), .B(B[14]), .Ci(\CTMP[14] ), .S(S[14]), .Co(
        \CTMP[15] ) );
  FA_174 FA_i_16 ( .A(A[15]), .B(B[15]), .Ci(\CTMP[15] ), .S(S[15]), .Co(
        \CTMP[16] ) );
  FA_173 FA_i_17 ( .A(A[16]), .B(B[16]), .Ci(\CTMP[16] ), .S(S[16]), .Co(
        \CTMP[17] ) );
  FA_172 FA_i_18 ( .A(A[17]), .B(B[17]), .Ci(\CTMP[17] ), .S(S[17]), .Co(
        \CTMP[18] ) );
  FA_171 FA_i_19 ( .A(A[18]), .B(B[18]), .Ci(\CTMP[18] ), .S(S[18]), .Co(
        \CTMP[19] ) );
  FA_170 FA_i_20 ( .A(A[19]), .B(B[19]), .Ci(\CTMP[19] ), .S(S[19]), .Co(
        \CTMP[20] ) );
  FA_169 FA_i_21 ( .A(A[20]), .B(B[20]), .Ci(\CTMP[20] ), .S(S[20]), .Co(
        \CTMP[21] ) );
  FA_168 FA_i_22 ( .A(A[21]), .B(B[21]), .Ci(\CTMP[21] ), .S(S[21]), .Co(
        \CTMP[22] ) );
  FA_167 FA_i_23 ( .A(A[22]), .B(B[22]), .Ci(\CTMP[22] ), .S(S[22]), .Co(
        \CTMP[23] ) );
  FA_166 FA_i_24 ( .A(A[23]), .B(B[23]), .Ci(\CTMP[23] ), .S(S[23]), .Co(
        \CTMP[24] ) );
  FA_165 FA_i_25 ( .A(A[24]), .B(B[24]), .Ci(\CTMP[24] ), .S(S[24]), .Co(
        \CTMP[25] ) );
  FA_164 FA_i_26 ( .A(A[25]), .B(B[25]), .Ci(\CTMP[25] ), .S(S[25]), .Co(
        \CTMP[26] ) );
  FA_163 FA_i_27 ( .A(A[26]), .B(B[26]), .Ci(\CTMP[26] ), .S(S[26]), .Co(
        \CTMP[27] ) );
  FA_162 FA_i_28 ( .A(A[27]), .B(B[27]), .Ci(\CTMP[27] ), .S(S[27]), .Co(
        \CTMP[28] ) );
  FA_161 FA_i_29 ( .A(A[28]), .B(B[28]), .Ci(\CTMP[28] ), .S(S[28]), .Co(
        \CTMP[29] ) );
  FA_160 FA_i_30 ( .A(A[29]), .B(B[29]), .Ci(\CTMP[29] ), .S(S[29]), .Co(Co)
         );
endmodule


module mux5to1_N30 ( A, B, C, D, E, Y, SEL );
  input [29:0] A;
  input [29:0] B;
  input [29:0] C;
  input [29:0] D;
  input [29:0] E;
  output [29:0] Y;
  input [2:0] SEL;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299;

  BUF_X1 U1 ( .A(n8), .Z(n289) );
  BUF_X1 U2 ( .A(n8), .Z(n288) );
  BUF_X1 U3 ( .A(n9), .Z(n286) );
  BUF_X1 U4 ( .A(n9), .Z(n285) );
  BUF_X1 U5 ( .A(n6), .Z(n295) );
  BUF_X1 U6 ( .A(n6), .Z(n294) );
  BUF_X1 U7 ( .A(n7), .Z(n292) );
  BUF_X1 U8 ( .A(n7), .Z(n291) );
  BUF_X1 U9 ( .A(n5), .Z(n298) );
  BUF_X1 U10 ( .A(n5), .Z(n297) );
  BUF_X1 U11 ( .A(n9), .Z(n287) );
  BUF_X1 U12 ( .A(n8), .Z(n290) );
  BUF_X1 U13 ( .A(n6), .Z(n296) );
  BUF_X1 U14 ( .A(n7), .Z(n293) );
  BUF_X1 U15 ( .A(n5), .Z(n299) );
  NOR3_X1 U16 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n68), .ZN(n6) );
  NOR3_X1 U17 ( .A1(n68), .A2(SEL[2]), .A3(n69), .ZN(n7) );
  NOR3_X1 U18 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n69), .ZN(n8) );
  NOR2_X1 U19 ( .A1(n70), .A2(n287), .ZN(n5) );
  AOI21_X1 U20 ( .B1(n68), .B2(n69), .A(SEL[2]), .ZN(n70) );
  INV_X1 U21 ( .A(SEL[0]), .ZN(n69) );
  INV_X1 U22 ( .A(SEL[1]), .ZN(n68) );
  AND3_X1 U23 ( .A1(n69), .A2(n68), .A3(SEL[2]), .ZN(n9) );
  NAND2_X1 U24 ( .A1(n3), .A2(n4), .ZN(Y[9]) );
  AOI22_X1 U25 ( .A1(B[9]), .A2(n290), .B1(E[9]), .B2(n286), .ZN(n3) );
  AOI222_X1 U26 ( .A1(A[9]), .A2(n299), .B1(C[9]), .B2(n296), .C1(D[9]), .C2(
        n293), .ZN(n4) );
  NAND2_X1 U27 ( .A1(n10), .A2(n11), .ZN(Y[8]) );
  AOI22_X1 U28 ( .A1(B[8]), .A2(n290), .B1(E[8]), .B2(n285), .ZN(n10) );
  AOI222_X1 U29 ( .A1(A[8]), .A2(n299), .B1(C[8]), .B2(n296), .C1(D[8]), .C2(
        n293), .ZN(n11) );
  NAND2_X1 U30 ( .A1(n12), .A2(n13), .ZN(Y[7]) );
  AOI22_X1 U31 ( .A1(B[7]), .A2(n290), .B1(E[7]), .B2(n285), .ZN(n12) );
  AOI222_X1 U32 ( .A1(A[7]), .A2(n299), .B1(C[7]), .B2(n296), .C1(D[7]), .C2(
        n293), .ZN(n13) );
  NAND2_X1 U33 ( .A1(n14), .A2(n15), .ZN(Y[6]) );
  AOI22_X1 U34 ( .A1(B[6]), .A2(n290), .B1(E[6]), .B2(n285), .ZN(n14) );
  AOI222_X1 U35 ( .A1(A[6]), .A2(n299), .B1(C[6]), .B2(n296), .C1(D[6]), .C2(
        n293), .ZN(n15) );
  NAND2_X1 U36 ( .A1(n16), .A2(n17), .ZN(Y[5]) );
  AOI22_X1 U37 ( .A1(B[5]), .A2(n290), .B1(E[5]), .B2(n285), .ZN(n16) );
  AOI222_X1 U38 ( .A1(A[5]), .A2(n299), .B1(C[5]), .B2(n296), .C1(D[5]), .C2(
        n293), .ZN(n17) );
  NAND2_X1 U39 ( .A1(n18), .A2(n19), .ZN(Y[4]) );
  AOI22_X1 U40 ( .A1(B[4]), .A2(n290), .B1(E[4]), .B2(n285), .ZN(n18) );
  AOI222_X1 U41 ( .A1(A[4]), .A2(n299), .B1(C[4]), .B2(n296), .C1(D[4]), .C2(
        n293), .ZN(n19) );
  NAND2_X1 U42 ( .A1(n24), .A2(n25), .ZN(Y[29]) );
  AOI22_X1 U43 ( .A1(B[29]), .A2(n289), .B1(E[29]), .B2(n285), .ZN(n24) );
  AOI222_X1 U44 ( .A1(A[29]), .A2(n298), .B1(C[29]), .B2(n295), .C1(D[29]), 
        .C2(n292), .ZN(n25) );
  NAND2_X1 U45 ( .A1(n26), .A2(n27), .ZN(Y[28]) );
  AOI22_X1 U46 ( .A1(B[28]), .A2(n289), .B1(E[28]), .B2(n285), .ZN(n26) );
  AOI222_X1 U47 ( .A1(A[28]), .A2(n298), .B1(C[28]), .B2(n295), .C1(D[28]), 
        .C2(n292), .ZN(n27) );
  NAND2_X1 U48 ( .A1(n28), .A2(n29), .ZN(Y[27]) );
  AOI22_X1 U49 ( .A1(B[27]), .A2(n289), .B1(E[27]), .B2(n285), .ZN(n28) );
  AOI222_X1 U50 ( .A1(A[27]), .A2(n298), .B1(C[27]), .B2(n295), .C1(D[27]), 
        .C2(n292), .ZN(n29) );
  NAND2_X1 U51 ( .A1(n30), .A2(n31), .ZN(Y[26]) );
  AOI22_X1 U52 ( .A1(B[26]), .A2(n289), .B1(E[26]), .B2(n285), .ZN(n30) );
  AOI222_X1 U53 ( .A1(A[26]), .A2(n298), .B1(C[26]), .B2(n295), .C1(D[26]), 
        .C2(n292), .ZN(n31) );
  NAND2_X1 U54 ( .A1(n32), .A2(n33), .ZN(Y[25]) );
  AOI22_X1 U55 ( .A1(B[25]), .A2(n289), .B1(E[25]), .B2(n286), .ZN(n32) );
  AOI222_X1 U56 ( .A1(A[25]), .A2(n298), .B1(C[25]), .B2(n295), .C1(D[25]), 
        .C2(n292), .ZN(n33) );
  NAND2_X1 U57 ( .A1(n34), .A2(n35), .ZN(Y[24]) );
  AOI22_X1 U58 ( .A1(B[24]), .A2(n289), .B1(E[24]), .B2(n286), .ZN(n34) );
  AOI222_X1 U59 ( .A1(A[24]), .A2(n298), .B1(C[24]), .B2(n295), .C1(D[24]), 
        .C2(n292), .ZN(n35) );
  NAND2_X1 U60 ( .A1(n36), .A2(n37), .ZN(Y[23]) );
  AOI22_X1 U61 ( .A1(B[23]), .A2(n289), .B1(E[23]), .B2(n286), .ZN(n36) );
  AOI222_X1 U62 ( .A1(A[23]), .A2(n298), .B1(C[23]), .B2(n295), .C1(D[23]), 
        .C2(n292), .ZN(n37) );
  NAND2_X1 U63 ( .A1(n38), .A2(n39), .ZN(Y[22]) );
  AOI22_X1 U64 ( .A1(B[22]), .A2(n289), .B1(E[22]), .B2(n286), .ZN(n38) );
  AOI222_X1 U65 ( .A1(A[22]), .A2(n298), .B1(C[22]), .B2(n295), .C1(D[22]), 
        .C2(n292), .ZN(n39) );
  NAND2_X1 U66 ( .A1(n40), .A2(n41), .ZN(Y[21]) );
  AOI22_X1 U67 ( .A1(B[21]), .A2(n289), .B1(E[21]), .B2(n286), .ZN(n40) );
  AOI222_X1 U68 ( .A1(A[21]), .A2(n298), .B1(C[21]), .B2(n295), .C1(D[21]), 
        .C2(n292), .ZN(n41) );
  NAND2_X1 U69 ( .A1(n42), .A2(n43), .ZN(Y[20]) );
  AOI22_X1 U70 ( .A1(B[20]), .A2(n289), .B1(E[20]), .B2(n286), .ZN(n42) );
  AOI222_X1 U71 ( .A1(A[20]), .A2(n298), .B1(C[20]), .B2(n295), .C1(D[20]), 
        .C2(n292), .ZN(n43) );
  NAND2_X1 U72 ( .A1(n46), .A2(n47), .ZN(Y[19]) );
  AOI22_X1 U73 ( .A1(B[19]), .A2(n288), .B1(E[19]), .B2(n286), .ZN(n46) );
  AOI222_X1 U74 ( .A1(A[19]), .A2(n297), .B1(C[19]), .B2(n294), .C1(D[19]), 
        .C2(n291), .ZN(n47) );
  NAND2_X1 U75 ( .A1(n48), .A2(n49), .ZN(Y[18]) );
  AOI22_X1 U76 ( .A1(B[18]), .A2(n288), .B1(E[18]), .B2(n286), .ZN(n48) );
  AOI222_X1 U77 ( .A1(A[18]), .A2(n297), .B1(C[18]), .B2(n294), .C1(D[18]), 
        .C2(n291), .ZN(n49) );
  NAND2_X1 U78 ( .A1(n50), .A2(n51), .ZN(Y[17]) );
  AOI22_X1 U79 ( .A1(B[17]), .A2(n288), .B1(E[17]), .B2(n286), .ZN(n50) );
  AOI222_X1 U80 ( .A1(A[17]), .A2(n297), .B1(C[17]), .B2(n294), .C1(D[17]), 
        .C2(n291), .ZN(n51) );
  NAND2_X1 U81 ( .A1(n52), .A2(n53), .ZN(Y[16]) );
  AOI22_X1 U82 ( .A1(B[16]), .A2(n288), .B1(E[16]), .B2(n286), .ZN(n52) );
  AOI222_X1 U83 ( .A1(A[16]), .A2(n297), .B1(C[16]), .B2(n294), .C1(D[16]), 
        .C2(n291), .ZN(n53) );
  NAND2_X1 U84 ( .A1(n54), .A2(n55), .ZN(Y[15]) );
  AOI22_X1 U85 ( .A1(B[15]), .A2(n288), .B1(E[15]), .B2(n287), .ZN(n54) );
  AOI222_X1 U86 ( .A1(A[15]), .A2(n297), .B1(C[15]), .B2(n294), .C1(D[15]), 
        .C2(n291), .ZN(n55) );
  NAND2_X1 U87 ( .A1(n56), .A2(n57), .ZN(Y[14]) );
  AOI22_X1 U88 ( .A1(B[14]), .A2(n288), .B1(E[14]), .B2(n287), .ZN(n56) );
  AOI222_X1 U89 ( .A1(A[14]), .A2(n297), .B1(C[14]), .B2(n294), .C1(D[14]), 
        .C2(n291), .ZN(n57) );
  NAND2_X1 U90 ( .A1(n58), .A2(n59), .ZN(Y[13]) );
  AOI22_X1 U91 ( .A1(B[13]), .A2(n288), .B1(E[13]), .B2(n287), .ZN(n58) );
  AOI222_X1 U92 ( .A1(A[13]), .A2(n297), .B1(C[13]), .B2(n294), .C1(D[13]), 
        .C2(n291), .ZN(n59) );
  NAND2_X1 U93 ( .A1(n60), .A2(n61), .ZN(Y[12]) );
  AOI22_X1 U94 ( .A1(B[12]), .A2(n288), .B1(E[12]), .B2(n287), .ZN(n60) );
  AOI222_X1 U95 ( .A1(A[12]), .A2(n297), .B1(C[12]), .B2(n294), .C1(D[12]), 
        .C2(n291), .ZN(n61) );
  NAND2_X1 U96 ( .A1(n62), .A2(n63), .ZN(Y[11]) );
  AOI22_X1 U97 ( .A1(B[11]), .A2(n288), .B1(E[11]), .B2(n287), .ZN(n62) );
  AOI222_X1 U98 ( .A1(A[11]), .A2(n297), .B1(C[11]), .B2(n294), .C1(D[11]), 
        .C2(n291), .ZN(n63) );
  NAND2_X1 U99 ( .A1(n64), .A2(n65), .ZN(Y[10]) );
  AOI22_X1 U100 ( .A1(B[10]), .A2(n288), .B1(E[10]), .B2(n287), .ZN(n64) );
  AOI222_X1 U101 ( .A1(A[10]), .A2(n297), .B1(C[10]), .B2(n294), .C1(D[10]), 
        .C2(n291), .ZN(n65) );
  NAND2_X1 U102 ( .A1(n20), .A2(n21), .ZN(Y[3]) );
  AOI22_X1 U103 ( .A1(B[3]), .A2(n289), .B1(E[3]), .B2(n285), .ZN(n20) );
  AOI222_X1 U104 ( .A1(A[3]), .A2(n298), .B1(C[3]), .B2(n295), .C1(D[3]), .C2(
        n292), .ZN(n21) );
  NAND2_X1 U105 ( .A1(n22), .A2(n23), .ZN(Y[2]) );
  AOI22_X1 U106 ( .A1(B[2]), .A2(n289), .B1(E[2]), .B2(n285), .ZN(n22) );
  AOI222_X1 U107 ( .A1(A[2]), .A2(n298), .B1(C[2]), .B2(n295), .C1(D[2]), .C2(
        n292), .ZN(n23) );
  NAND2_X1 U108 ( .A1(n44), .A2(n45), .ZN(Y[1]) );
  AOI22_X1 U109 ( .A1(B[1]), .A2(n288), .B1(E[1]), .B2(n286), .ZN(n44) );
  AOI222_X1 U110 ( .A1(A[1]), .A2(n297), .B1(C[1]), .B2(n294), .C1(D[1]), .C2(
        n291), .ZN(n45) );
  NAND2_X1 U111 ( .A1(n66), .A2(n67), .ZN(Y[0]) );
  AOI22_X1 U112 ( .A1(B[0]), .A2(n288), .B1(E[0]), .B2(n285), .ZN(n66) );
  AOI222_X1 U113 ( .A1(A[0]), .A2(n297), .B1(C[0]), .B2(n294), .C1(D[0]), .C2(
        n291), .ZN(n67) );
endmodule


module rca_N28 ( A, B, S, Co );
  input [27:0] A;
  input [27:0] B;
  output [27:0] S;
  output Co;
  wire   \CTMP[9] , \CTMP[8] , \CTMP[7] , \CTMP[6] , \CTMP[5] , \CTMP[4] ,
         \CTMP[3] , \CTMP[2] , \CTMP[27] , \CTMP[26] , \CTMP[25] , \CTMP[24] ,
         \CTMP[23] , \CTMP[22] , \CTMP[21] , \CTMP[20] , \CTMP[1] , \CTMP[19] ,
         \CTMP[18] , \CTMP[17] , \CTMP[16] , \CTMP[15] , \CTMP[14] ,
         \CTMP[13] , \CTMP[12] , \CTMP[11] , \CTMP[10] ;

  HA_3 HA_0 ( .A(A[0]), .B(B[0]), .S(S[0]), .Co(\CTMP[1] ) );
  FA_215 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(\CTMP[1] ), .S(S[1]), .Co(\CTMP[2] )
         );
  FA_214 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(\CTMP[2] ), .S(S[2]), .Co(\CTMP[3] )
         );
  FA_213 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(\CTMP[3] ), .S(S[3]), .Co(\CTMP[4] )
         );
  FA_212 FA_i_5 ( .A(A[4]), .B(B[4]), .Ci(\CTMP[4] ), .S(S[4]), .Co(\CTMP[5] )
         );
  FA_211 FA_i_6 ( .A(A[5]), .B(B[5]), .Ci(\CTMP[5] ), .S(S[5]), .Co(\CTMP[6] )
         );
  FA_210 FA_i_7 ( .A(A[6]), .B(B[6]), .Ci(\CTMP[6] ), .S(S[6]), .Co(\CTMP[7] )
         );
  FA_209 FA_i_8 ( .A(A[7]), .B(B[7]), .Ci(\CTMP[7] ), .S(S[7]), .Co(\CTMP[8] )
         );
  FA_208 FA_i_9 ( .A(A[8]), .B(B[8]), .Ci(\CTMP[8] ), .S(S[8]), .Co(\CTMP[9] )
         );
  FA_207 FA_i_10 ( .A(A[9]), .B(B[9]), .Ci(\CTMP[9] ), .S(S[9]), .Co(
        \CTMP[10] ) );
  FA_206 FA_i_11 ( .A(A[10]), .B(B[10]), .Ci(\CTMP[10] ), .S(S[10]), .Co(
        \CTMP[11] ) );
  FA_205 FA_i_12 ( .A(A[11]), .B(B[11]), .Ci(\CTMP[11] ), .S(S[11]), .Co(
        \CTMP[12] ) );
  FA_204 FA_i_13 ( .A(A[12]), .B(B[12]), .Ci(\CTMP[12] ), .S(S[12]), .Co(
        \CTMP[13] ) );
  FA_203 FA_i_14 ( .A(A[13]), .B(B[13]), .Ci(\CTMP[13] ), .S(S[13]), .Co(
        \CTMP[14] ) );
  FA_202 FA_i_15 ( .A(A[14]), .B(B[14]), .Ci(\CTMP[14] ), .S(S[14]), .Co(
        \CTMP[15] ) );
  FA_201 FA_i_16 ( .A(A[15]), .B(B[15]), .Ci(\CTMP[15] ), .S(S[15]), .Co(
        \CTMP[16] ) );
  FA_200 FA_i_17 ( .A(A[16]), .B(B[16]), .Ci(\CTMP[16] ), .S(S[16]), .Co(
        \CTMP[17] ) );
  FA_199 FA_i_18 ( .A(A[17]), .B(B[17]), .Ci(\CTMP[17] ), .S(S[17]), .Co(
        \CTMP[18] ) );
  FA_198 FA_i_19 ( .A(A[18]), .B(B[18]), .Ci(\CTMP[18] ), .S(S[18]), .Co(
        \CTMP[19] ) );
  FA_197 FA_i_20 ( .A(A[19]), .B(B[19]), .Ci(\CTMP[19] ), .S(S[19]), .Co(
        \CTMP[20] ) );
  FA_196 FA_i_21 ( .A(A[20]), .B(B[20]), .Ci(\CTMP[20] ), .S(S[20]), .Co(
        \CTMP[21] ) );
  FA_195 FA_i_22 ( .A(A[21]), .B(B[21]), .Ci(\CTMP[21] ), .S(S[21]), .Co(
        \CTMP[22] ) );
  FA_194 FA_i_23 ( .A(A[22]), .B(B[22]), .Ci(\CTMP[22] ), .S(S[22]), .Co(
        \CTMP[23] ) );
  FA_193 FA_i_24 ( .A(A[23]), .B(B[23]), .Ci(\CTMP[23] ), .S(S[23]), .Co(
        \CTMP[24] ) );
  FA_192 FA_i_25 ( .A(A[24]), .B(B[24]), .Ci(\CTMP[24] ), .S(S[24]), .Co(
        \CTMP[25] ) );
  FA_191 FA_i_26 ( .A(A[25]), .B(B[25]), .Ci(\CTMP[25] ), .S(S[25]), .Co(
        \CTMP[26] ) );
  FA_190 FA_i_27 ( .A(A[26]), .B(B[26]), .Ci(\CTMP[26] ), .S(S[26]), .Co(
        \CTMP[27] ) );
  FA_189 FA_i_28 ( .A(A[27]), .B(B[27]), .Ci(\CTMP[27] ), .S(S[27]), .Co(Co)
         );
endmodule


module mux5to1_N28 ( A, B, C, D, E, Y, SEL );
  input [27:0] A;
  input [27:0] B;
  input [27:0] C;
  input [27:0] D;
  input [27:0] E;
  output [27:0] Y;
  input [2:0] SEL;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287;

  BUF_X1 U1 ( .A(n8), .Z(n277) );
  BUF_X1 U2 ( .A(n8), .Z(n276) );
  BUF_X1 U3 ( .A(n9), .Z(n273) );
  BUF_X1 U4 ( .A(n9), .Z(n274) );
  BUF_X1 U5 ( .A(n6), .Z(n283) );
  BUF_X1 U6 ( .A(n6), .Z(n282) );
  BUF_X1 U7 ( .A(n7), .Z(n280) );
  BUF_X1 U8 ( .A(n7), .Z(n279) );
  BUF_X1 U9 ( .A(n5), .Z(n286) );
  BUF_X1 U10 ( .A(n5), .Z(n285) );
  BUF_X1 U11 ( .A(n9), .Z(n275) );
  BUF_X1 U12 ( .A(n8), .Z(n278) );
  BUF_X1 U13 ( .A(n6), .Z(n284) );
  BUF_X1 U14 ( .A(n7), .Z(n281) );
  BUF_X1 U15 ( .A(n5), .Z(n287) );
  NOR3_X1 U16 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n64), .ZN(n6) );
  NOR3_X1 U17 ( .A1(n64), .A2(SEL[2]), .A3(n65), .ZN(n7) );
  NOR3_X1 U18 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n65), .ZN(n8) );
  NOR2_X1 U19 ( .A1(n66), .A2(n275), .ZN(n5) );
  AOI21_X1 U20 ( .B1(n64), .B2(n65), .A(SEL[2]), .ZN(n66) );
  INV_X1 U21 ( .A(SEL[0]), .ZN(n65) );
  INV_X1 U22 ( .A(SEL[1]), .ZN(n64) );
  AND3_X1 U23 ( .A1(n65), .A2(n64), .A3(SEL[2]), .ZN(n9) );
  NAND2_X1 U24 ( .A1(n24), .A2(n25), .ZN(Y[27]) );
  AOI22_X1 U25 ( .A1(B[27]), .A2(n277), .B1(E[27]), .B2(n274), .ZN(n24) );
  AOI222_X1 U26 ( .A1(A[27]), .A2(n286), .B1(C[27]), .B2(n283), .C1(D[27]), 
        .C2(n280), .ZN(n25) );
  NAND2_X1 U27 ( .A1(n26), .A2(n27), .ZN(Y[26]) );
  AOI22_X1 U28 ( .A1(B[26]), .A2(n277), .B1(E[26]), .B2(n274), .ZN(n26) );
  AOI222_X1 U29 ( .A1(A[26]), .A2(n286), .B1(C[26]), .B2(n283), .C1(D[26]), 
        .C2(n280), .ZN(n27) );
  NAND2_X1 U30 ( .A1(n28), .A2(n29), .ZN(Y[25]) );
  AOI22_X1 U31 ( .A1(B[25]), .A2(n277), .B1(E[25]), .B2(n274), .ZN(n28) );
  AOI222_X1 U32 ( .A1(A[25]), .A2(n286), .B1(C[25]), .B2(n283), .C1(D[25]), 
        .C2(n280), .ZN(n29) );
  NAND2_X1 U33 ( .A1(n30), .A2(n31), .ZN(Y[24]) );
  AOI22_X1 U34 ( .A1(B[24]), .A2(n277), .B1(E[24]), .B2(n274), .ZN(n30) );
  AOI222_X1 U35 ( .A1(A[24]), .A2(n286), .B1(C[24]), .B2(n283), .C1(D[24]), 
        .C2(n280), .ZN(n31) );
  NAND2_X1 U36 ( .A1(n32), .A2(n33), .ZN(Y[23]) );
  AOI22_X1 U37 ( .A1(B[23]), .A2(n277), .B1(E[23]), .B2(n274), .ZN(n32) );
  AOI222_X1 U38 ( .A1(A[23]), .A2(n286), .B1(C[23]), .B2(n283), .C1(D[23]), 
        .C2(n280), .ZN(n33) );
  NAND2_X1 U39 ( .A1(n34), .A2(n35), .ZN(Y[22]) );
  AOI22_X1 U40 ( .A1(B[22]), .A2(n277), .B1(E[22]), .B2(n274), .ZN(n34) );
  AOI222_X1 U41 ( .A1(A[22]), .A2(n286), .B1(C[22]), .B2(n283), .C1(D[22]), 
        .C2(n280), .ZN(n35) );
  NAND2_X1 U42 ( .A1(n36), .A2(n37), .ZN(Y[21]) );
  AOI22_X1 U43 ( .A1(B[21]), .A2(n277), .B1(E[21]), .B2(n274), .ZN(n36) );
  AOI222_X1 U44 ( .A1(A[21]), .A2(n286), .B1(C[21]), .B2(n283), .C1(D[21]), 
        .C2(n280), .ZN(n37) );
  NAND2_X1 U45 ( .A1(n38), .A2(n39), .ZN(Y[20]) );
  AOI22_X1 U46 ( .A1(B[20]), .A2(n277), .B1(E[20]), .B2(n274), .ZN(n38) );
  AOI222_X1 U47 ( .A1(A[20]), .A2(n286), .B1(C[20]), .B2(n283), .C1(D[20]), 
        .C2(n280), .ZN(n39) );
  NAND2_X1 U48 ( .A1(n42), .A2(n43), .ZN(Y[19]) );
  AOI22_X1 U49 ( .A1(B[19]), .A2(n276), .B1(E[19]), .B2(n273), .ZN(n42) );
  AOI222_X1 U50 ( .A1(A[19]), .A2(n285), .B1(C[19]), .B2(n282), .C1(D[19]), 
        .C2(n279), .ZN(n43) );
  NAND2_X1 U51 ( .A1(n44), .A2(n45), .ZN(Y[18]) );
  AOI22_X1 U52 ( .A1(B[18]), .A2(n276), .B1(E[18]), .B2(n273), .ZN(n44) );
  AOI222_X1 U53 ( .A1(A[18]), .A2(n285), .B1(C[18]), .B2(n282), .C1(D[18]), 
        .C2(n279), .ZN(n45) );
  NAND2_X1 U54 ( .A1(n46), .A2(n47), .ZN(Y[17]) );
  AOI22_X1 U55 ( .A1(B[17]), .A2(n276), .B1(E[17]), .B2(n273), .ZN(n46) );
  AOI222_X1 U56 ( .A1(A[17]), .A2(n285), .B1(C[17]), .B2(n282), .C1(D[17]), 
        .C2(n279), .ZN(n47) );
  NAND2_X1 U57 ( .A1(n48), .A2(n49), .ZN(Y[16]) );
  AOI22_X1 U58 ( .A1(B[16]), .A2(n276), .B1(E[16]), .B2(n273), .ZN(n48) );
  AOI222_X1 U59 ( .A1(A[16]), .A2(n285), .B1(C[16]), .B2(n282), .C1(D[16]), 
        .C2(n279), .ZN(n49) );
  NAND2_X1 U60 ( .A1(n50), .A2(n51), .ZN(Y[15]) );
  AOI22_X1 U61 ( .A1(B[15]), .A2(n276), .B1(E[15]), .B2(n273), .ZN(n50) );
  AOI222_X1 U62 ( .A1(A[15]), .A2(n285), .B1(C[15]), .B2(n282), .C1(D[15]), 
        .C2(n279), .ZN(n51) );
  NAND2_X1 U63 ( .A1(n52), .A2(n53), .ZN(Y[14]) );
  AOI22_X1 U64 ( .A1(B[14]), .A2(n276), .B1(E[14]), .B2(n273), .ZN(n52) );
  AOI222_X1 U65 ( .A1(A[14]), .A2(n285), .B1(C[14]), .B2(n282), .C1(D[14]), 
        .C2(n279), .ZN(n53) );
  NAND2_X1 U66 ( .A1(n54), .A2(n55), .ZN(Y[13]) );
  AOI22_X1 U67 ( .A1(B[13]), .A2(n276), .B1(E[13]), .B2(n273), .ZN(n54) );
  AOI222_X1 U68 ( .A1(A[13]), .A2(n285), .B1(C[13]), .B2(n282), .C1(D[13]), 
        .C2(n279), .ZN(n55) );
  NAND2_X1 U69 ( .A1(n56), .A2(n57), .ZN(Y[12]) );
  AOI22_X1 U70 ( .A1(B[12]), .A2(n276), .B1(E[12]), .B2(n273), .ZN(n56) );
  AOI222_X1 U71 ( .A1(A[12]), .A2(n285), .B1(C[12]), .B2(n282), .C1(D[12]), 
        .C2(n279), .ZN(n57) );
  NAND2_X1 U72 ( .A1(n58), .A2(n59), .ZN(Y[11]) );
  AOI22_X1 U73 ( .A1(B[11]), .A2(n276), .B1(E[11]), .B2(n273), .ZN(n58) );
  AOI222_X1 U74 ( .A1(A[11]), .A2(n285), .B1(C[11]), .B2(n282), .C1(D[11]), 
        .C2(n279), .ZN(n59) );
  NAND2_X1 U75 ( .A1(n60), .A2(n61), .ZN(Y[10]) );
  AOI22_X1 U76 ( .A1(B[10]), .A2(n276), .B1(E[10]), .B2(n273), .ZN(n60) );
  AOI222_X1 U77 ( .A1(A[10]), .A2(n285), .B1(C[10]), .B2(n282), .C1(D[10]), 
        .C2(n279), .ZN(n61) );
  NAND2_X1 U78 ( .A1(n3), .A2(n4), .ZN(Y[9]) );
  AOI22_X1 U79 ( .A1(B[9]), .A2(n278), .B1(E[9]), .B2(n273), .ZN(n3) );
  AOI222_X1 U80 ( .A1(A[9]), .A2(n287), .B1(C[9]), .B2(n284), .C1(D[9]), .C2(
        n281), .ZN(n4) );
  NAND2_X1 U81 ( .A1(n10), .A2(n11), .ZN(Y[8]) );
  AOI22_X1 U82 ( .A1(B[8]), .A2(n278), .B1(E[8]), .B2(n275), .ZN(n10) );
  AOI222_X1 U83 ( .A1(A[8]), .A2(n287), .B1(C[8]), .B2(n284), .C1(D[8]), .C2(
        n281), .ZN(n11) );
  NAND2_X1 U84 ( .A1(n12), .A2(n13), .ZN(Y[7]) );
  AOI22_X1 U85 ( .A1(B[7]), .A2(n278), .B1(E[7]), .B2(n275), .ZN(n12) );
  AOI222_X1 U86 ( .A1(A[7]), .A2(n287), .B1(C[7]), .B2(n284), .C1(D[7]), .C2(
        n281), .ZN(n13) );
  NAND2_X1 U87 ( .A1(n14), .A2(n15), .ZN(Y[6]) );
  AOI22_X1 U88 ( .A1(B[6]), .A2(n278), .B1(E[6]), .B2(n275), .ZN(n14) );
  AOI222_X1 U89 ( .A1(A[6]), .A2(n287), .B1(C[6]), .B2(n284), .C1(D[6]), .C2(
        n281), .ZN(n15) );
  NAND2_X1 U90 ( .A1(n16), .A2(n17), .ZN(Y[5]) );
  AOI22_X1 U91 ( .A1(B[5]), .A2(n277), .B1(E[5]), .B2(n275), .ZN(n16) );
  AOI222_X1 U92 ( .A1(A[5]), .A2(n286), .B1(C[5]), .B2(n283), .C1(D[5]), .C2(
        n280), .ZN(n17) );
  NAND2_X1 U93 ( .A1(n18), .A2(n19), .ZN(Y[4]) );
  AOI22_X1 U94 ( .A1(B[4]), .A2(n277), .B1(E[4]), .B2(n274), .ZN(n18) );
  AOI222_X1 U95 ( .A1(A[4]), .A2(n286), .B1(C[4]), .B2(n283), .C1(D[4]), .C2(
        n280), .ZN(n19) );
  NAND2_X1 U96 ( .A1(n20), .A2(n21), .ZN(Y[3]) );
  AOI22_X1 U97 ( .A1(B[3]), .A2(n277), .B1(E[3]), .B2(n274), .ZN(n20) );
  AOI222_X1 U98 ( .A1(A[3]), .A2(n286), .B1(C[3]), .B2(n283), .C1(D[3]), .C2(
        n280), .ZN(n21) );
  NAND2_X1 U99 ( .A1(n22), .A2(n23), .ZN(Y[2]) );
  AOI22_X1 U100 ( .A1(B[2]), .A2(n277), .B1(E[2]), .B2(n274), .ZN(n22) );
  AOI222_X1 U101 ( .A1(A[2]), .A2(n286), .B1(C[2]), .B2(n283), .C1(D[2]), .C2(
        n280), .ZN(n23) );
  NAND2_X1 U102 ( .A1(n40), .A2(n41), .ZN(Y[1]) );
  AOI22_X1 U103 ( .A1(B[1]), .A2(n276), .B1(E[1]), .B2(n273), .ZN(n40) );
  AOI222_X1 U104 ( .A1(A[1]), .A2(n285), .B1(C[1]), .B2(n282), .C1(D[1]), .C2(
        n279), .ZN(n41) );
  NAND2_X1 U105 ( .A1(n62), .A2(n63), .ZN(Y[0]) );
  AOI22_X1 U106 ( .A1(B[0]), .A2(n276), .B1(E[0]), .B2(n274), .ZN(n62) );
  AOI222_X1 U107 ( .A1(A[0]), .A2(n285), .B1(C[0]), .B2(n282), .C1(D[0]), .C2(
        n279), .ZN(n63) );
endmodule


module rca_N26 ( A, B, S, Co );
  input [25:0] A;
  input [25:0] B;
  output [25:0] S;
  output Co;
  wire   \CTMP[9] , \CTMP[8] , \CTMP[7] , \CTMP[6] , \CTMP[5] , \CTMP[4] ,
         \CTMP[3] , \CTMP[2] , \CTMP[25] , \CTMP[24] , \CTMP[23] , \CTMP[22] ,
         \CTMP[21] , \CTMP[20] , \CTMP[1] , \CTMP[19] , \CTMP[18] , \CTMP[17] ,
         \CTMP[16] , \CTMP[15] , \CTMP[14] , \CTMP[13] , \CTMP[12] ,
         \CTMP[11] , \CTMP[10] ;

  HA_4 HA_0 ( .A(A[0]), .B(B[0]), .S(S[0]), .Co(\CTMP[1] ) );
  FA_240 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(\CTMP[1] ), .S(S[1]), .Co(\CTMP[2] )
         );
  FA_239 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(\CTMP[2] ), .S(S[2]), .Co(\CTMP[3] )
         );
  FA_238 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(\CTMP[3] ), .S(S[3]), .Co(\CTMP[4] )
         );
  FA_237 FA_i_5 ( .A(A[4]), .B(B[4]), .Ci(\CTMP[4] ), .S(S[4]), .Co(\CTMP[5] )
         );
  FA_236 FA_i_6 ( .A(A[5]), .B(B[5]), .Ci(\CTMP[5] ), .S(S[5]), .Co(\CTMP[6] )
         );
  FA_235 FA_i_7 ( .A(A[6]), .B(B[6]), .Ci(\CTMP[6] ), .S(S[6]), .Co(\CTMP[7] )
         );
  FA_234 FA_i_8 ( .A(A[7]), .B(B[7]), .Ci(\CTMP[7] ), .S(S[7]), .Co(\CTMP[8] )
         );
  FA_233 FA_i_9 ( .A(A[8]), .B(B[8]), .Ci(\CTMP[8] ), .S(S[8]), .Co(\CTMP[9] )
         );
  FA_232 FA_i_10 ( .A(A[9]), .B(B[9]), .Ci(\CTMP[9] ), .S(S[9]), .Co(
        \CTMP[10] ) );
  FA_231 FA_i_11 ( .A(A[10]), .B(B[10]), .Ci(\CTMP[10] ), .S(S[10]), .Co(
        \CTMP[11] ) );
  FA_230 FA_i_12 ( .A(A[11]), .B(B[11]), .Ci(\CTMP[11] ), .S(S[11]), .Co(
        \CTMP[12] ) );
  FA_229 FA_i_13 ( .A(A[12]), .B(B[12]), .Ci(\CTMP[12] ), .S(S[12]), .Co(
        \CTMP[13] ) );
  FA_228 FA_i_14 ( .A(A[13]), .B(B[13]), .Ci(\CTMP[13] ), .S(S[13]), .Co(
        \CTMP[14] ) );
  FA_227 FA_i_15 ( .A(A[14]), .B(B[14]), .Ci(\CTMP[14] ), .S(S[14]), .Co(
        \CTMP[15] ) );
  FA_226 FA_i_16 ( .A(A[15]), .B(B[15]), .Ci(\CTMP[15] ), .S(S[15]), .Co(
        \CTMP[16] ) );
  FA_225 FA_i_17 ( .A(A[16]), .B(B[16]), .Ci(\CTMP[16] ), .S(S[16]), .Co(
        \CTMP[17] ) );
  FA_224 FA_i_18 ( .A(A[17]), .B(B[17]), .Ci(\CTMP[17] ), .S(S[17]), .Co(
        \CTMP[18] ) );
  FA_223 FA_i_19 ( .A(A[18]), .B(B[18]), .Ci(\CTMP[18] ), .S(S[18]), .Co(
        \CTMP[19] ) );
  FA_222 FA_i_20 ( .A(A[19]), .B(B[19]), .Ci(\CTMP[19] ), .S(S[19]), .Co(
        \CTMP[20] ) );
  FA_221 FA_i_21 ( .A(A[20]), .B(B[20]), .Ci(\CTMP[20] ), .S(S[20]), .Co(
        \CTMP[21] ) );
  FA_220 FA_i_22 ( .A(A[21]), .B(B[21]), .Ci(\CTMP[21] ), .S(S[21]), .Co(
        \CTMP[22] ) );
  FA_219 FA_i_23 ( .A(A[22]), .B(B[22]), .Ci(\CTMP[22] ), .S(S[22]), .Co(
        \CTMP[23] ) );
  FA_218 FA_i_24 ( .A(A[23]), .B(B[23]), .Ci(\CTMP[23] ), .S(S[23]), .Co(
        \CTMP[24] ) );
  FA_217 FA_i_25 ( .A(A[24]), .B(B[24]), .Ci(\CTMP[24] ), .S(S[24]), .Co(
        \CTMP[25] ) );
  FA_216 FA_i_26 ( .A(A[25]), .B(B[25]), .Ci(\CTMP[25] ), .S(S[25]), .Co(Co)
         );
endmodule


module mux5to1_N26 ( A, B, C, D, E, Y, SEL );
  input [25:0] A;
  input [25:0] B;
  input [25:0] C;
  input [25:0] D;
  input [25:0] E;
  output [25:0] Y;
  input [2:0] SEL;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271;

  BUF_X1 U1 ( .A(n8), .Z(n261) );
  BUF_X1 U2 ( .A(n8), .Z(n260) );
  BUF_X1 U3 ( .A(n9), .Z(n257) );
  BUF_X1 U4 ( .A(n9), .Z(n258) );
  BUF_X1 U5 ( .A(n6), .Z(n267) );
  BUF_X1 U6 ( .A(n6), .Z(n266) );
  BUF_X1 U7 ( .A(n7), .Z(n264) );
  BUF_X1 U8 ( .A(n7), .Z(n263) );
  BUF_X1 U9 ( .A(n5), .Z(n270) );
  BUF_X1 U10 ( .A(n5), .Z(n269) );
  BUF_X1 U11 ( .A(n9), .Z(n259) );
  BUF_X1 U12 ( .A(n8), .Z(n262) );
  BUF_X1 U13 ( .A(n6), .Z(n268) );
  BUF_X1 U14 ( .A(n7), .Z(n265) );
  BUF_X1 U15 ( .A(n5), .Z(n271) );
  NOR3_X1 U16 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n60), .ZN(n6) );
  NOR3_X1 U17 ( .A1(n60), .A2(SEL[2]), .A3(n61), .ZN(n7) );
  NOR3_X1 U18 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n61), .ZN(n8) );
  NOR2_X1 U19 ( .A1(n62), .A2(n259), .ZN(n5) );
  AOI21_X1 U20 ( .B1(n60), .B2(n61), .A(SEL[2]), .ZN(n62) );
  INV_X1 U21 ( .A(SEL[0]), .ZN(n61) );
  INV_X1 U22 ( .A(SEL[1]), .ZN(n60) );
  AND3_X1 U23 ( .A1(n61), .A2(n60), .A3(SEL[2]), .ZN(n9) );
  NAND2_X1 U24 ( .A1(n24), .A2(n25), .ZN(Y[25]) );
  AOI22_X1 U25 ( .A1(B[25]), .A2(n261), .B1(E[25]), .B2(n258), .ZN(n24) );
  AOI222_X1 U26 ( .A1(A[25]), .A2(n270), .B1(C[25]), .B2(n267), .C1(D[25]), 
        .C2(n264), .ZN(n25) );
  NAND2_X1 U27 ( .A1(n26), .A2(n27), .ZN(Y[24]) );
  AOI22_X1 U28 ( .A1(B[24]), .A2(n261), .B1(E[24]), .B2(n258), .ZN(n26) );
  AOI222_X1 U29 ( .A1(A[24]), .A2(n270), .B1(C[24]), .B2(n267), .C1(D[24]), 
        .C2(n264), .ZN(n27) );
  NAND2_X1 U30 ( .A1(n28), .A2(n29), .ZN(Y[23]) );
  AOI22_X1 U31 ( .A1(B[23]), .A2(n261), .B1(E[23]), .B2(n258), .ZN(n28) );
  AOI222_X1 U32 ( .A1(A[23]), .A2(n270), .B1(C[23]), .B2(n267), .C1(D[23]), 
        .C2(n264), .ZN(n29) );
  NAND2_X1 U33 ( .A1(n30), .A2(n31), .ZN(Y[22]) );
  AOI22_X1 U34 ( .A1(B[22]), .A2(n261), .B1(E[22]), .B2(n258), .ZN(n30) );
  AOI222_X1 U35 ( .A1(A[22]), .A2(n270), .B1(C[22]), .B2(n267), .C1(D[22]), 
        .C2(n264), .ZN(n31) );
  NAND2_X1 U36 ( .A1(n32), .A2(n33), .ZN(Y[21]) );
  AOI22_X1 U37 ( .A1(B[21]), .A2(n261), .B1(E[21]), .B2(n258), .ZN(n32) );
  AOI222_X1 U38 ( .A1(A[21]), .A2(n270), .B1(C[21]), .B2(n267), .C1(D[21]), 
        .C2(n264), .ZN(n33) );
  NAND2_X1 U39 ( .A1(n34), .A2(n35), .ZN(Y[20]) );
  AOI22_X1 U40 ( .A1(B[20]), .A2(n261), .B1(E[20]), .B2(n258), .ZN(n34) );
  AOI222_X1 U41 ( .A1(A[20]), .A2(n270), .B1(C[20]), .B2(n267), .C1(D[20]), 
        .C2(n264), .ZN(n35) );
  NAND2_X1 U42 ( .A1(n38), .A2(n39), .ZN(Y[19]) );
  AOI22_X1 U43 ( .A1(B[19]), .A2(n260), .B1(E[19]), .B2(n257), .ZN(n38) );
  AOI222_X1 U44 ( .A1(A[19]), .A2(n269), .B1(C[19]), .B2(n266), .C1(D[19]), 
        .C2(n263), .ZN(n39) );
  NAND2_X1 U45 ( .A1(n40), .A2(n41), .ZN(Y[18]) );
  AOI22_X1 U46 ( .A1(B[18]), .A2(n260), .B1(E[18]), .B2(n257), .ZN(n40) );
  AOI222_X1 U47 ( .A1(A[18]), .A2(n269), .B1(C[18]), .B2(n266), .C1(D[18]), 
        .C2(n263), .ZN(n41) );
  NAND2_X1 U48 ( .A1(n42), .A2(n43), .ZN(Y[17]) );
  AOI22_X1 U49 ( .A1(B[17]), .A2(n260), .B1(E[17]), .B2(n257), .ZN(n42) );
  AOI222_X1 U50 ( .A1(A[17]), .A2(n269), .B1(C[17]), .B2(n266), .C1(D[17]), 
        .C2(n263), .ZN(n43) );
  NAND2_X1 U51 ( .A1(n44), .A2(n45), .ZN(Y[16]) );
  AOI22_X1 U52 ( .A1(B[16]), .A2(n260), .B1(E[16]), .B2(n257), .ZN(n44) );
  AOI222_X1 U53 ( .A1(A[16]), .A2(n269), .B1(C[16]), .B2(n266), .C1(D[16]), 
        .C2(n263), .ZN(n45) );
  NAND2_X1 U54 ( .A1(n46), .A2(n47), .ZN(Y[15]) );
  AOI22_X1 U55 ( .A1(B[15]), .A2(n260), .B1(E[15]), .B2(n257), .ZN(n46) );
  AOI222_X1 U56 ( .A1(A[15]), .A2(n269), .B1(C[15]), .B2(n266), .C1(D[15]), 
        .C2(n263), .ZN(n47) );
  NAND2_X1 U57 ( .A1(n48), .A2(n49), .ZN(Y[14]) );
  AOI22_X1 U58 ( .A1(B[14]), .A2(n260), .B1(E[14]), .B2(n257), .ZN(n48) );
  AOI222_X1 U59 ( .A1(A[14]), .A2(n269), .B1(C[14]), .B2(n266), .C1(D[14]), 
        .C2(n263), .ZN(n49) );
  NAND2_X1 U60 ( .A1(n50), .A2(n51), .ZN(Y[13]) );
  AOI22_X1 U61 ( .A1(B[13]), .A2(n260), .B1(E[13]), .B2(n257), .ZN(n50) );
  AOI222_X1 U62 ( .A1(A[13]), .A2(n269), .B1(C[13]), .B2(n266), .C1(D[13]), 
        .C2(n263), .ZN(n51) );
  NAND2_X1 U63 ( .A1(n52), .A2(n53), .ZN(Y[12]) );
  AOI22_X1 U64 ( .A1(B[12]), .A2(n260), .B1(E[12]), .B2(n257), .ZN(n52) );
  AOI222_X1 U65 ( .A1(A[12]), .A2(n269), .B1(C[12]), .B2(n266), .C1(D[12]), 
        .C2(n263), .ZN(n53) );
  NAND2_X1 U66 ( .A1(n54), .A2(n55), .ZN(Y[11]) );
  AOI22_X1 U67 ( .A1(B[11]), .A2(n260), .B1(E[11]), .B2(n257), .ZN(n54) );
  AOI222_X1 U68 ( .A1(A[11]), .A2(n269), .B1(C[11]), .B2(n266), .C1(D[11]), 
        .C2(n263), .ZN(n55) );
  NAND2_X1 U69 ( .A1(n56), .A2(n57), .ZN(Y[10]) );
  AOI22_X1 U70 ( .A1(B[10]), .A2(n260), .B1(E[10]), .B2(n257), .ZN(n56) );
  AOI222_X1 U71 ( .A1(A[10]), .A2(n269), .B1(C[10]), .B2(n266), .C1(D[10]), 
        .C2(n263), .ZN(n57) );
  NAND2_X1 U72 ( .A1(n12), .A2(n13), .ZN(Y[7]) );
  AOI22_X1 U73 ( .A1(B[7]), .A2(n261), .B1(E[7]), .B2(n259), .ZN(n12) );
  AOI222_X1 U74 ( .A1(A[7]), .A2(n270), .B1(C[7]), .B2(n267), .C1(D[7]), .C2(
        n264), .ZN(n13) );
  NAND2_X1 U75 ( .A1(n14), .A2(n15), .ZN(Y[6]) );
  AOI22_X1 U76 ( .A1(B[6]), .A2(n261), .B1(E[6]), .B2(n258), .ZN(n14) );
  AOI222_X1 U77 ( .A1(A[6]), .A2(n270), .B1(C[6]), .B2(n267), .C1(D[6]), .C2(
        n264), .ZN(n15) );
  NAND2_X1 U78 ( .A1(n16), .A2(n17), .ZN(Y[5]) );
  AOI22_X1 U79 ( .A1(B[5]), .A2(n261), .B1(E[5]), .B2(n258), .ZN(n16) );
  AOI222_X1 U80 ( .A1(A[5]), .A2(n270), .B1(C[5]), .B2(n267), .C1(D[5]), .C2(
        n264), .ZN(n17) );
  NAND2_X1 U81 ( .A1(n18), .A2(n19), .ZN(Y[4]) );
  AOI22_X1 U82 ( .A1(B[4]), .A2(n261), .B1(E[4]), .B2(n258), .ZN(n18) );
  AOI222_X1 U83 ( .A1(A[4]), .A2(n270), .B1(C[4]), .B2(n267), .C1(D[4]), .C2(
        n264), .ZN(n19) );
  NAND2_X1 U84 ( .A1(n20), .A2(n21), .ZN(Y[3]) );
  AOI22_X1 U85 ( .A1(B[3]), .A2(n261), .B1(E[3]), .B2(n258), .ZN(n20) );
  AOI222_X1 U86 ( .A1(A[3]), .A2(n270), .B1(C[3]), .B2(n267), .C1(D[3]), .C2(
        n264), .ZN(n21) );
  NAND2_X1 U87 ( .A1(n22), .A2(n23), .ZN(Y[2]) );
  AOI22_X1 U88 ( .A1(B[2]), .A2(n261), .B1(E[2]), .B2(n258), .ZN(n22) );
  AOI222_X1 U89 ( .A1(A[2]), .A2(n270), .B1(C[2]), .B2(n267), .C1(D[2]), .C2(
        n264), .ZN(n23) );
  NAND2_X1 U90 ( .A1(n36), .A2(n37), .ZN(Y[1]) );
  AOI22_X1 U91 ( .A1(B[1]), .A2(n260), .B1(E[1]), .B2(n257), .ZN(n36) );
  AOI222_X1 U92 ( .A1(A[1]), .A2(n269), .B1(C[1]), .B2(n266), .C1(D[1]), .C2(
        n263), .ZN(n37) );
  NAND2_X1 U93 ( .A1(n58), .A2(n59), .ZN(Y[0]) );
  AOI22_X1 U94 ( .A1(B[0]), .A2(n260), .B1(E[0]), .B2(n258), .ZN(n58) );
  AOI222_X1 U95 ( .A1(A[0]), .A2(n269), .B1(C[0]), .B2(n266), .C1(D[0]), .C2(
        n263), .ZN(n59) );
  NAND2_X1 U96 ( .A1(n3), .A2(n4), .ZN(Y[9]) );
  AOI22_X1 U97 ( .A1(B[9]), .A2(n262), .B1(E[9]), .B2(n257), .ZN(n3) );
  AOI222_X1 U98 ( .A1(A[9]), .A2(n271), .B1(C[9]), .B2(n268), .C1(D[9]), .C2(
        n265), .ZN(n4) );
  NAND2_X1 U99 ( .A1(n10), .A2(n11), .ZN(Y[8]) );
  AOI22_X1 U100 ( .A1(B[8]), .A2(n262), .B1(E[8]), .B2(n259), .ZN(n10) );
  AOI222_X1 U101 ( .A1(A[8]), .A2(n271), .B1(C[8]), .B2(n268), .C1(D[8]), .C2(
        n265), .ZN(n11) );
endmodule


module rca_N24 ( A, B, S, Co );
  input [23:0] A;
  input [23:0] B;
  output [23:0] S;
  output Co;
  wire   \CTMP[9] , \CTMP[8] , \CTMP[7] , \CTMP[6] , \CTMP[5] , \CTMP[4] ,
         \CTMP[3] , \CTMP[2] , \CTMP[23] , \CTMP[22] , \CTMP[21] , \CTMP[20] ,
         \CTMP[1] , \CTMP[19] , \CTMP[18] , \CTMP[17] , \CTMP[16] , \CTMP[15] ,
         \CTMP[14] , \CTMP[13] , \CTMP[12] , \CTMP[11] , \CTMP[10] ;

  HA_5 HA_0 ( .A(A[0]), .B(B[0]), .S(S[0]), .Co(\CTMP[1] ) );
  FA_263 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(\CTMP[1] ), .S(S[1]), .Co(\CTMP[2] )
         );
  FA_262 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(\CTMP[2] ), .S(S[2]), .Co(\CTMP[3] )
         );
  FA_261 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(\CTMP[3] ), .S(S[3]), .Co(\CTMP[4] )
         );
  FA_260 FA_i_5 ( .A(A[4]), .B(B[4]), .Ci(\CTMP[4] ), .S(S[4]), .Co(\CTMP[5] )
         );
  FA_259 FA_i_6 ( .A(A[5]), .B(B[5]), .Ci(\CTMP[5] ), .S(S[5]), .Co(\CTMP[6] )
         );
  FA_258 FA_i_7 ( .A(A[6]), .B(B[6]), .Ci(\CTMP[6] ), .S(S[6]), .Co(\CTMP[7] )
         );
  FA_257 FA_i_8 ( .A(A[7]), .B(B[7]), .Ci(\CTMP[7] ), .S(S[7]), .Co(\CTMP[8] )
         );
  FA_256 FA_i_9 ( .A(A[8]), .B(B[8]), .Ci(\CTMP[8] ), .S(S[8]), .Co(\CTMP[9] )
         );
  FA_255 FA_i_10 ( .A(A[9]), .B(B[9]), .Ci(\CTMP[9] ), .S(S[9]), .Co(
        \CTMP[10] ) );
  FA_254 FA_i_11 ( .A(A[10]), .B(B[10]), .Ci(\CTMP[10] ), .S(S[10]), .Co(
        \CTMP[11] ) );
  FA_253 FA_i_12 ( .A(A[11]), .B(B[11]), .Ci(\CTMP[11] ), .S(S[11]), .Co(
        \CTMP[12] ) );
  FA_252 FA_i_13 ( .A(A[12]), .B(B[12]), .Ci(\CTMP[12] ), .S(S[12]), .Co(
        \CTMP[13] ) );
  FA_251 FA_i_14 ( .A(A[13]), .B(B[13]), .Ci(\CTMP[13] ), .S(S[13]), .Co(
        \CTMP[14] ) );
  FA_250 FA_i_15 ( .A(A[14]), .B(B[14]), .Ci(\CTMP[14] ), .S(S[14]), .Co(
        \CTMP[15] ) );
  FA_249 FA_i_16 ( .A(A[15]), .B(B[15]), .Ci(\CTMP[15] ), .S(S[15]), .Co(
        \CTMP[16] ) );
  FA_248 FA_i_17 ( .A(A[16]), .B(B[16]), .Ci(\CTMP[16] ), .S(S[16]), .Co(
        \CTMP[17] ) );
  FA_247 FA_i_18 ( .A(A[17]), .B(B[17]), .Ci(\CTMP[17] ), .S(S[17]), .Co(
        \CTMP[18] ) );
  FA_246 FA_i_19 ( .A(A[18]), .B(B[18]), .Ci(\CTMP[18] ), .S(S[18]), .Co(
        \CTMP[19] ) );
  FA_245 FA_i_20 ( .A(A[19]), .B(B[19]), .Ci(\CTMP[19] ), .S(S[19]), .Co(
        \CTMP[20] ) );
  FA_244 FA_i_21 ( .A(A[20]), .B(B[20]), .Ci(\CTMP[20] ), .S(S[20]), .Co(
        \CTMP[21] ) );
  FA_243 FA_i_22 ( .A(A[21]), .B(B[21]), .Ci(\CTMP[21] ), .S(S[21]), .Co(
        \CTMP[22] ) );
  FA_242 FA_i_23 ( .A(A[22]), .B(B[22]), .Ci(\CTMP[22] ), .S(S[22]), .Co(
        \CTMP[23] ) );
  FA_241 FA_i_24 ( .A(A[23]), .B(B[23]), .Ci(\CTMP[23] ), .S(S[23]), .Co(Co)
         );
endmodule


module mux5to1_N24 ( A, B, C, D, E, Y, SEL );
  input [23:0] A;
  input [23:0] B;
  input [23:0] C;
  input [23:0] D;
  input [23:0] E;
  output [23:0] Y;
  input [2:0] SEL;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172;

  BUF_X1 U1 ( .A(n7), .Z(n168) );
  BUF_X1 U2 ( .A(n7), .Z(n167) );
  BUF_X1 U3 ( .A(n8), .Z(n166) );
  BUF_X1 U4 ( .A(n8), .Z(n165) );
  BUF_X1 U5 ( .A(n9), .Z(n164) );
  BUF_X1 U6 ( .A(n9), .Z(n163) );
  BUF_X1 U7 ( .A(n6), .Z(n170) );
  BUF_X1 U8 ( .A(n6), .Z(n169) );
  BUF_X1 U9 ( .A(n5), .Z(n171) );
  BUF_X1 U10 ( .A(n5), .Z(n172) );
  NOR3_X1 U11 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n58), .ZN(n8) );
  NOR3_X1 U12 ( .A1(n56), .A2(SEL[2]), .A3(n58), .ZN(n9) );
  NOR3_X1 U13 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n56), .ZN(n7) );
  NOR2_X1 U14 ( .A1(n57), .A2(n171), .ZN(n6) );
  AOI21_X1 U15 ( .B1(n58), .B2(n56), .A(SEL[2]), .ZN(n57) );
  INV_X1 U16 ( .A(SEL[0]), .ZN(n56) );
  INV_X1 U17 ( .A(SEL[1]), .ZN(n58) );
  AND3_X1 U18 ( .A1(n56), .A2(n58), .A3(SEL[2]), .ZN(n5) );
  NAND2_X1 U19 ( .A1(n24), .A2(n25), .ZN(Y[23]) );
  AOI22_X1 U20 ( .A1(C[23]), .A2(n166), .B1(D[23]), .B2(n164), .ZN(n24) );
  AOI222_X1 U21 ( .A1(E[23]), .A2(n172), .B1(A[23]), .B2(n170), .C1(B[23]), 
        .C2(n168), .ZN(n25) );
  NAND2_X1 U22 ( .A1(n26), .A2(n27), .ZN(Y[22]) );
  AOI22_X1 U23 ( .A1(C[22]), .A2(n166), .B1(D[22]), .B2(n164), .ZN(n26) );
  AOI222_X1 U24 ( .A1(E[22]), .A2(n172), .B1(A[22]), .B2(n170), .C1(B[22]), 
        .C2(n168), .ZN(n27) );
  NAND2_X1 U25 ( .A1(n28), .A2(n29), .ZN(Y[21]) );
  AOI22_X1 U26 ( .A1(C[21]), .A2(n166), .B1(D[21]), .B2(n164), .ZN(n28) );
  AOI222_X1 U27 ( .A1(E[21]), .A2(n172), .B1(A[21]), .B2(n170), .C1(B[21]), 
        .C2(n168), .ZN(n29) );
  NAND2_X1 U28 ( .A1(n30), .A2(n31), .ZN(Y[20]) );
  AOI22_X1 U29 ( .A1(C[20]), .A2(n166), .B1(D[20]), .B2(n164), .ZN(n30) );
  AOI222_X1 U30 ( .A1(E[20]), .A2(n172), .B1(A[20]), .B2(n170), .C1(B[20]), 
        .C2(n168), .ZN(n31) );
  NAND2_X1 U31 ( .A1(n34), .A2(n35), .ZN(Y[19]) );
  AOI22_X1 U32 ( .A1(C[19]), .A2(n165), .B1(D[19]), .B2(n163), .ZN(n34) );
  AOI222_X1 U33 ( .A1(E[19]), .A2(n171), .B1(A[19]), .B2(n169), .C1(B[19]), 
        .C2(n167), .ZN(n35) );
  NAND2_X1 U34 ( .A1(n36), .A2(n37), .ZN(Y[18]) );
  AOI22_X1 U35 ( .A1(C[18]), .A2(n165), .B1(D[18]), .B2(n163), .ZN(n36) );
  AOI222_X1 U36 ( .A1(E[18]), .A2(n171), .B1(A[18]), .B2(n169), .C1(B[18]), 
        .C2(n167), .ZN(n37) );
  NAND2_X1 U37 ( .A1(n38), .A2(n39), .ZN(Y[17]) );
  AOI22_X1 U38 ( .A1(C[17]), .A2(n165), .B1(D[17]), .B2(n163), .ZN(n38) );
  AOI222_X1 U39 ( .A1(E[17]), .A2(n171), .B1(A[17]), .B2(n169), .C1(B[17]), 
        .C2(n167), .ZN(n39) );
  NAND2_X1 U40 ( .A1(n40), .A2(n41), .ZN(Y[16]) );
  AOI22_X1 U41 ( .A1(C[16]), .A2(n165), .B1(D[16]), .B2(n163), .ZN(n40) );
  AOI222_X1 U42 ( .A1(E[16]), .A2(n171), .B1(A[16]), .B2(n169), .C1(B[16]), 
        .C2(n167), .ZN(n41) );
  NAND2_X1 U43 ( .A1(n42), .A2(n43), .ZN(Y[15]) );
  AOI22_X1 U44 ( .A1(C[15]), .A2(n165), .B1(D[15]), .B2(n163), .ZN(n42) );
  AOI222_X1 U45 ( .A1(E[15]), .A2(n171), .B1(A[15]), .B2(n169), .C1(B[15]), 
        .C2(n167), .ZN(n43) );
  NAND2_X1 U46 ( .A1(n44), .A2(n45), .ZN(Y[14]) );
  AOI22_X1 U47 ( .A1(C[14]), .A2(n165), .B1(D[14]), .B2(n163), .ZN(n44) );
  AOI222_X1 U48 ( .A1(E[14]), .A2(n171), .B1(A[14]), .B2(n169), .C1(B[14]), 
        .C2(n167), .ZN(n45) );
  NAND2_X1 U49 ( .A1(n46), .A2(n47), .ZN(Y[13]) );
  AOI22_X1 U50 ( .A1(C[13]), .A2(n165), .B1(D[13]), .B2(n163), .ZN(n46) );
  AOI222_X1 U51 ( .A1(E[13]), .A2(n171), .B1(A[13]), .B2(n169), .C1(B[13]), 
        .C2(n167), .ZN(n47) );
  NAND2_X1 U52 ( .A1(n48), .A2(n49), .ZN(Y[12]) );
  AOI22_X1 U53 ( .A1(C[12]), .A2(n165), .B1(D[12]), .B2(n163), .ZN(n48) );
  AOI222_X1 U54 ( .A1(E[12]), .A2(n171), .B1(A[12]), .B2(n169), .C1(B[12]), 
        .C2(n167), .ZN(n49) );
  NAND2_X1 U55 ( .A1(n50), .A2(n51), .ZN(Y[11]) );
  AOI22_X1 U56 ( .A1(C[11]), .A2(n165), .B1(D[11]), .B2(n163), .ZN(n50) );
  AOI222_X1 U57 ( .A1(E[11]), .A2(n171), .B1(A[11]), .B2(n169), .C1(B[11]), 
        .C2(n167), .ZN(n51) );
  NAND2_X1 U58 ( .A1(n52), .A2(n53), .ZN(Y[10]) );
  AOI22_X1 U59 ( .A1(C[10]), .A2(n165), .B1(D[10]), .B2(n163), .ZN(n52) );
  AOI222_X1 U60 ( .A1(E[10]), .A2(n171), .B1(A[10]), .B2(n169), .C1(B[10]), 
        .C2(n167), .ZN(n53) );
  NAND2_X1 U61 ( .A1(n3), .A2(n4), .ZN(Y[9]) );
  AOI22_X1 U62 ( .A1(C[9]), .A2(n166), .B1(D[9]), .B2(n164), .ZN(n3) );
  AOI222_X1 U63 ( .A1(E[9]), .A2(n5), .B1(A[9]), .B2(n170), .C1(B[9]), .C2(
        n168), .ZN(n4) );
  NAND2_X1 U64 ( .A1(n10), .A2(n11), .ZN(Y[8]) );
  AOI22_X1 U65 ( .A1(C[8]), .A2(n166), .B1(D[8]), .B2(n164), .ZN(n10) );
  AOI222_X1 U66 ( .A1(E[8]), .A2(n172), .B1(A[8]), .B2(n170), .C1(B[8]), .C2(
        n168), .ZN(n11) );
  NAND2_X1 U67 ( .A1(n12), .A2(n13), .ZN(Y[7]) );
  AOI22_X1 U68 ( .A1(C[7]), .A2(n166), .B1(D[7]), .B2(n164), .ZN(n12) );
  AOI222_X1 U69 ( .A1(E[7]), .A2(n172), .B1(A[7]), .B2(n170), .C1(B[7]), .C2(
        n168), .ZN(n13) );
  NAND2_X1 U70 ( .A1(n14), .A2(n15), .ZN(Y[6]) );
  AOI22_X1 U71 ( .A1(C[6]), .A2(n166), .B1(D[6]), .B2(n164), .ZN(n14) );
  AOI222_X1 U72 ( .A1(E[6]), .A2(n172), .B1(A[6]), .B2(n170), .C1(B[6]), .C2(
        n168), .ZN(n15) );
  NAND2_X1 U73 ( .A1(n16), .A2(n17), .ZN(Y[5]) );
  AOI22_X1 U74 ( .A1(C[5]), .A2(n166), .B1(D[5]), .B2(n164), .ZN(n16) );
  AOI222_X1 U75 ( .A1(E[5]), .A2(n172), .B1(A[5]), .B2(n170), .C1(B[5]), .C2(
        n168), .ZN(n17) );
  NAND2_X1 U76 ( .A1(n18), .A2(n19), .ZN(Y[4]) );
  AOI22_X1 U77 ( .A1(C[4]), .A2(n166), .B1(D[4]), .B2(n164), .ZN(n18) );
  AOI222_X1 U78 ( .A1(E[4]), .A2(n172), .B1(A[4]), .B2(n170), .C1(B[4]), .C2(
        n168), .ZN(n19) );
  NAND2_X1 U79 ( .A1(n20), .A2(n21), .ZN(Y[3]) );
  AOI22_X1 U80 ( .A1(C[3]), .A2(n166), .B1(D[3]), .B2(n164), .ZN(n20) );
  AOI222_X1 U81 ( .A1(E[3]), .A2(n172), .B1(A[3]), .B2(n170), .C1(B[3]), .C2(
        n168), .ZN(n21) );
  NAND2_X1 U82 ( .A1(n22), .A2(n23), .ZN(Y[2]) );
  AOI22_X1 U83 ( .A1(C[2]), .A2(n166), .B1(D[2]), .B2(n164), .ZN(n22) );
  AOI222_X1 U84 ( .A1(E[2]), .A2(n172), .B1(A[2]), .B2(n170), .C1(B[2]), .C2(
        n168), .ZN(n23) );
  NAND2_X1 U85 ( .A1(n32), .A2(n33), .ZN(Y[1]) );
  AOI22_X1 U86 ( .A1(C[1]), .A2(n165), .B1(D[1]), .B2(n163), .ZN(n32) );
  AOI222_X1 U87 ( .A1(E[1]), .A2(n172), .B1(A[1]), .B2(n169), .C1(B[1]), .C2(
        n167), .ZN(n33) );
  NAND2_X1 U88 ( .A1(n54), .A2(n55), .ZN(Y[0]) );
  AOI22_X1 U89 ( .A1(C[0]), .A2(n165), .B1(D[0]), .B2(n163), .ZN(n54) );
  AOI222_X1 U90 ( .A1(E[0]), .A2(n171), .B1(A[0]), .B2(n169), .C1(B[0]), .C2(
        n167), .ZN(n55) );
endmodule


module rca_N22 ( A, B, S, Co );
  input [21:0] A;
  input [21:0] B;
  output [21:0] S;
  output Co;
  wire   \CTMP[9] , \CTMP[8] , \CTMP[7] , \CTMP[6] , \CTMP[5] , \CTMP[4] ,
         \CTMP[3] , \CTMP[2] , \CTMP[21] , \CTMP[20] , \CTMP[1] , \CTMP[19] ,
         \CTMP[18] , \CTMP[17] , \CTMP[16] , \CTMP[15] , \CTMP[14] ,
         \CTMP[13] , \CTMP[12] , \CTMP[11] , \CTMP[10] ;

  HA_6 HA_0 ( .A(A[0]), .B(B[0]), .S(S[0]), .Co(\CTMP[1] ) );
  FA_284 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(\CTMP[1] ), .S(S[1]), .Co(\CTMP[2] )
         );
  FA_283 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(\CTMP[2] ), .S(S[2]), .Co(\CTMP[3] )
         );
  FA_282 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(\CTMP[3] ), .S(S[3]), .Co(\CTMP[4] )
         );
  FA_281 FA_i_5 ( .A(A[4]), .B(B[4]), .Ci(\CTMP[4] ), .S(S[4]), .Co(\CTMP[5] )
         );
  FA_280 FA_i_6 ( .A(A[5]), .B(B[5]), .Ci(\CTMP[5] ), .S(S[5]), .Co(\CTMP[6] )
         );
  FA_279 FA_i_7 ( .A(A[6]), .B(B[6]), .Ci(\CTMP[6] ), .S(S[6]), .Co(\CTMP[7] )
         );
  FA_278 FA_i_8 ( .A(A[7]), .B(B[7]), .Ci(\CTMP[7] ), .S(S[7]), .Co(\CTMP[8] )
         );
  FA_277 FA_i_9 ( .A(A[8]), .B(B[8]), .Ci(\CTMP[8] ), .S(S[8]), .Co(\CTMP[9] )
         );
  FA_276 FA_i_10 ( .A(A[9]), .B(B[9]), .Ci(\CTMP[9] ), .S(S[9]), .Co(
        \CTMP[10] ) );
  FA_275 FA_i_11 ( .A(A[10]), .B(B[10]), .Ci(\CTMP[10] ), .S(S[10]), .Co(
        \CTMP[11] ) );
  FA_274 FA_i_12 ( .A(A[11]), .B(B[11]), .Ci(\CTMP[11] ), .S(S[11]), .Co(
        \CTMP[12] ) );
  FA_273 FA_i_13 ( .A(A[12]), .B(B[12]), .Ci(\CTMP[12] ), .S(S[12]), .Co(
        \CTMP[13] ) );
  FA_272 FA_i_14 ( .A(A[13]), .B(B[13]), .Ci(\CTMP[13] ), .S(S[13]), .Co(
        \CTMP[14] ) );
  FA_271 FA_i_15 ( .A(A[14]), .B(B[14]), .Ci(\CTMP[14] ), .S(S[14]), .Co(
        \CTMP[15] ) );
  FA_270 FA_i_16 ( .A(A[15]), .B(B[15]), .Ci(\CTMP[15] ), .S(S[15]), .Co(
        \CTMP[16] ) );
  FA_269 FA_i_17 ( .A(A[16]), .B(B[16]), .Ci(\CTMP[16] ), .S(S[16]), .Co(
        \CTMP[17] ) );
  FA_268 FA_i_18 ( .A(A[17]), .B(B[17]), .Ci(\CTMP[17] ), .S(S[17]), .Co(
        \CTMP[18] ) );
  FA_267 FA_i_19 ( .A(A[18]), .B(B[18]), .Ci(\CTMP[18] ), .S(S[18]), .Co(
        \CTMP[19] ) );
  FA_266 FA_i_20 ( .A(A[19]), .B(B[19]), .Ci(\CTMP[19] ), .S(S[19]), .Co(
        \CTMP[20] ) );
  FA_265 FA_i_21 ( .A(A[20]), .B(B[20]), .Ci(\CTMP[20] ), .S(S[20]), .Co(
        \CTMP[21] ) );
  FA_264 FA_i_22 ( .A(A[21]), .B(B[21]), .Ci(\CTMP[21] ), .S(S[21]), .Co(Co)
         );
endmodule


module mux5to1_N22 ( A, B, C, D, E, Y, SEL );
  input [21:0] A;
  input [21:0] B;
  input [21:0] C;
  input [21:0] D;
  input [21:0] E;
  output [21:0] Y;
  input [2:0] SEL;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438;

  BUF_X1 U1 ( .A(n8), .Z(n415) );
  BUF_X1 U2 ( .A(n8), .Z(n414) );
  BUF_X1 U3 ( .A(n424), .Z(n428) );
  BUF_X1 U4 ( .A(n424), .Z(n427) );
  BUF_X1 U5 ( .A(n423), .Z(n426) );
  BUF_X1 U6 ( .A(n423), .Z(n425) );
  BUF_X1 U7 ( .A(n432), .Z(n436) );
  BUF_X1 U8 ( .A(n432), .Z(n435) );
  BUF_X1 U9 ( .A(n431), .Z(n434) );
  BUF_X1 U10 ( .A(n431), .Z(n433) );
  BUF_X1 U11 ( .A(n8), .Z(n417) );
  BUF_X1 U12 ( .A(n8), .Z(n416) );
  BUF_X1 U13 ( .A(n6), .Z(n430) );
  BUF_X1 U14 ( .A(n6), .Z(n429) );
  BUF_X1 U15 ( .A(n7), .Z(n438) );
  BUF_X1 U16 ( .A(n7), .Z(n437) );
  INV_X1 U17 ( .A(SEL[0]), .ZN(n53) );
  INV_X1 U18 ( .A(SEL[1]), .ZN(n52) );
  NOR3_X1 U19 ( .A1(n53), .A2(SEL[2]), .A3(n52), .ZN(n424) );
  NOR3_X1 U20 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n52), .ZN(n432) );
  NOR3_X1 U21 ( .A1(n53), .A2(SEL[2]), .A3(n52), .ZN(n6) );
  NOR3_X1 U22 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n52), .ZN(n7) );
  NOR3_X1 U23 ( .A1(n53), .A2(SEL[2]), .A3(n52), .ZN(n423) );
  NOR3_X1 U24 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n52), .ZN(n431) );
  NOR2_X1 U25 ( .A1(n54), .A2(n413), .ZN(n8) );
  AOI21_X1 U26 ( .B1(n52), .B2(n53), .A(SEL[2]), .ZN(n54) );
  BUF_X1 U27 ( .A(n418), .Z(n420) );
  NOR3_X1 U28 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n53), .ZN(n418) );
  BUF_X1 U29 ( .A(n419), .Z(n421) );
  NOR3_X1 U30 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n53), .ZN(n419) );
  BUF_X1 U31 ( .A(n5), .Z(n422) );
  NOR3_X1 U32 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n53), .ZN(n5) );
  AND3_X1 U33 ( .A1(n53), .A2(n52), .A3(SEL[2]), .ZN(n9) );
  NAND2_X1 U34 ( .A1(n24), .A2(n25), .ZN(Y[21]) );
  AOI22_X1 U35 ( .A1(A[21]), .A2(n417), .B1(E[21]), .B2(n406), .ZN(n24) );
  AOI222_X1 U36 ( .A1(B[21]), .A2(n421), .B1(D[21]), .B2(n428), .C1(C[21]), 
        .C2(n436), .ZN(n25) );
  NAND2_X1 U37 ( .A1(n26), .A2(n27), .ZN(Y[20]) );
  AOI22_X1 U38 ( .A1(A[20]), .A2(n416), .B1(E[20]), .B2(n407), .ZN(n26) );
  AOI222_X1 U39 ( .A1(B[20]), .A2(n421), .B1(D[20]), .B2(n427), .C1(C[20]), 
        .C2(n435), .ZN(n27) );
  NAND2_X1 U40 ( .A1(n30), .A2(n31), .ZN(Y[19]) );
  AOI22_X1 U41 ( .A1(A[19]), .A2(n414), .B1(E[19]), .B2(n408), .ZN(n30) );
  AOI222_X1 U42 ( .A1(B[19]), .A2(n422), .B1(D[19]), .B2(n425), .C1(C[19]), 
        .C2(n433), .ZN(n31) );
  NAND2_X1 U43 ( .A1(n32), .A2(n33), .ZN(Y[18]) );
  AOI22_X1 U44 ( .A1(A[18]), .A2(n415), .B1(E[18]), .B2(n413), .ZN(n32) );
  AOI222_X1 U45 ( .A1(B[18]), .A2(n420), .B1(D[18]), .B2(n426), .C1(C[18]), 
        .C2(n434), .ZN(n33) );
  NAND2_X1 U46 ( .A1(n34), .A2(n35), .ZN(Y[17]) );
  AOI22_X1 U47 ( .A1(A[17]), .A2(n414), .B1(E[17]), .B2(n409), .ZN(n34) );
  AOI222_X1 U48 ( .A1(B[17]), .A2(n421), .B1(D[17]), .B2(n425), .C1(C[17]), 
        .C2(n433), .ZN(n35) );
  NAND2_X1 U49 ( .A1(n36), .A2(n37), .ZN(Y[16]) );
  AOI22_X1 U50 ( .A1(A[16]), .A2(n417), .B1(E[16]), .B2(n412), .ZN(n36) );
  AOI222_X1 U51 ( .A1(B[16]), .A2(n420), .B1(D[16]), .B2(n430), .C1(C[16]), 
        .C2(n438), .ZN(n37) );
  NAND2_X1 U52 ( .A1(n38), .A2(n39), .ZN(Y[15]) );
  AOI22_X1 U53 ( .A1(A[15]), .A2(n416), .B1(E[15]), .B2(n411), .ZN(n38) );
  AOI222_X1 U54 ( .A1(B[15]), .A2(n422), .B1(D[15]), .B2(n429), .C1(C[15]), 
        .C2(n437), .ZN(n39) );
  NAND2_X1 U55 ( .A1(n40), .A2(n41), .ZN(Y[14]) );
  AOI22_X1 U56 ( .A1(A[14]), .A2(n417), .B1(E[14]), .B2(n411), .ZN(n40) );
  AOI222_X1 U57 ( .A1(B[14]), .A2(n422), .B1(D[14]), .B2(n430), .C1(C[14]), 
        .C2(n438), .ZN(n41) );
  NAND2_X1 U58 ( .A1(n42), .A2(n43), .ZN(Y[13]) );
  AOI22_X1 U59 ( .A1(A[13]), .A2(n416), .B1(E[13]), .B2(n410), .ZN(n42) );
  AOI222_X1 U60 ( .A1(B[13]), .A2(n421), .B1(D[13]), .B2(n429), .C1(C[13]), 
        .C2(n437), .ZN(n43) );
  NAND2_X1 U61 ( .A1(n44), .A2(n45), .ZN(Y[12]) );
  AOI22_X1 U62 ( .A1(A[12]), .A2(n415), .B1(E[12]), .B2(n409), .ZN(n44) );
  AOI222_X1 U63 ( .A1(B[12]), .A2(n421), .B1(D[12]), .B2(n428), .C1(C[12]), 
        .C2(n436), .ZN(n45) );
  NAND2_X1 U64 ( .A1(n46), .A2(n47), .ZN(Y[11]) );
  AOI22_X1 U65 ( .A1(A[11]), .A2(n414), .B1(E[11]), .B2(n408), .ZN(n46) );
  AOI222_X1 U66 ( .A1(B[11]), .A2(n420), .B1(D[11]), .B2(n427), .C1(C[11]), 
        .C2(n435), .ZN(n47) );
  NAND2_X1 U67 ( .A1(n48), .A2(n49), .ZN(Y[10]) );
  AOI22_X1 U68 ( .A1(A[10]), .A2(n415), .B1(E[10]), .B2(n407), .ZN(n48) );
  AOI222_X1 U69 ( .A1(B[10]), .A2(n422), .B1(D[10]), .B2(n426), .C1(C[10]), 
        .C2(n434), .ZN(n49) );
  NAND2_X1 U70 ( .A1(n3), .A2(n4), .ZN(Y[9]) );
  AOI22_X1 U71 ( .A1(A[9]), .A2(n417), .B1(E[9]), .B2(n412), .ZN(n3) );
  AOI222_X1 U72 ( .A1(B[9]), .A2(n421), .B1(D[9]), .B2(n428), .C1(C[9]), .C2(
        n436), .ZN(n4) );
  NAND2_X1 U73 ( .A1(n10), .A2(n11), .ZN(Y[8]) );
  AOI22_X1 U74 ( .A1(A[8]), .A2(n416), .B1(E[8]), .B2(n412), .ZN(n10) );
  AOI222_X1 U75 ( .A1(B[8]), .A2(n420), .B1(D[8]), .B2(n427), .C1(C[8]), .C2(
        n435), .ZN(n11) );
  NAND2_X1 U76 ( .A1(n12), .A2(n13), .ZN(Y[7]) );
  AOI22_X1 U77 ( .A1(A[7]), .A2(n415), .B1(E[7]), .B2(n411), .ZN(n12) );
  AOI222_X1 U78 ( .A1(B[7]), .A2(n422), .B1(D[7]), .B2(n426), .C1(C[7]), .C2(
        n434), .ZN(n13) );
  NAND2_X1 U79 ( .A1(n14), .A2(n15), .ZN(Y[6]) );
  AOI22_X1 U80 ( .A1(A[6]), .A2(n414), .B1(E[6]), .B2(n410), .ZN(n14) );
  AOI222_X1 U81 ( .A1(B[6]), .A2(n420), .B1(D[6]), .B2(n425), .C1(C[6]), .C2(
        n433), .ZN(n15) );
  NAND2_X1 U82 ( .A1(n16), .A2(n17), .ZN(Y[5]) );
  AOI22_X1 U83 ( .A1(A[5]), .A2(n415), .B1(E[5]), .B2(n409), .ZN(n16) );
  AOI222_X1 U84 ( .A1(B[5]), .A2(n421), .B1(D[5]), .B2(n428), .C1(C[5]), .C2(
        n436), .ZN(n17) );
  NAND2_X1 U85 ( .A1(n18), .A2(n19), .ZN(Y[4]) );
  AOI22_X1 U86 ( .A1(A[4]), .A2(n414), .B1(E[4]), .B2(n408), .ZN(n18) );
  AOI222_X1 U87 ( .A1(B[4]), .A2(n420), .B1(D[4]), .B2(n427), .C1(C[4]), .C2(
        n435), .ZN(n19) );
  NAND2_X1 U88 ( .A1(n20), .A2(n21), .ZN(Y[3]) );
  AOI22_X1 U89 ( .A1(A[3]), .A2(n417), .B1(E[3]), .B2(n407), .ZN(n20) );
  AOI222_X1 U90 ( .A1(B[3]), .A2(n422), .B1(D[3]), .B2(n430), .C1(C[3]), .C2(
        n438), .ZN(n21) );
  NAND2_X1 U91 ( .A1(n22), .A2(n23), .ZN(Y[2]) );
  AOI22_X1 U92 ( .A1(A[2]), .A2(n416), .B1(E[2]), .B2(n406), .ZN(n22) );
  AOI222_X1 U93 ( .A1(B[2]), .A2(n422), .B1(D[2]), .B2(n429), .C1(C[2]), .C2(
        n437), .ZN(n23) );
  NAND2_X1 U94 ( .A1(n28), .A2(n29), .ZN(Y[1]) );
  AOI22_X1 U95 ( .A1(A[1]), .A2(n415), .B1(E[1]), .B2(n410), .ZN(n28) );
  AOI222_X1 U96 ( .A1(B[1]), .A2(n420), .B1(D[1]), .B2(n426), .C1(C[1]), .C2(
        n434), .ZN(n29) );
  NAND2_X1 U97 ( .A1(n50), .A2(n51), .ZN(Y[0]) );
  AOI22_X1 U98 ( .A1(A[0]), .A2(n414), .B1(E[0]), .B2(n406), .ZN(n50) );
  AOI222_X1 U99 ( .A1(B[0]), .A2(n420), .B1(D[0]), .B2(n425), .C1(C[0]), .C2(
        n433), .ZN(n51) );
  INV_X1 U100 ( .A(n9), .ZN(n403) );
  INV_X1 U101 ( .A(n9), .ZN(n404) );
  INV_X1 U102 ( .A(n9), .ZN(n405) );
  INV_X1 U103 ( .A(n403), .ZN(n406) );
  INV_X1 U104 ( .A(n403), .ZN(n407) );
  INV_X1 U105 ( .A(n403), .ZN(n408) );
  INV_X1 U106 ( .A(n404), .ZN(n409) );
  INV_X1 U107 ( .A(n404), .ZN(n410) );
  INV_X1 U108 ( .A(n404), .ZN(n411) );
  INV_X1 U109 ( .A(n405), .ZN(n412) );
  INV_X1 U110 ( .A(n404), .ZN(n413) );
endmodule


module rca_N20 ( A, B, S, Co );
  input [19:0] A;
  input [19:0] B;
  output [19:0] S;
  output Co;
  wire   \CTMP[9] , \CTMP[8] , \CTMP[7] , \CTMP[6] , \CTMP[5] , \CTMP[4] ,
         \CTMP[3] , \CTMP[2] , \CTMP[1] , \CTMP[19] , \CTMP[18] , \CTMP[17] ,
         \CTMP[16] , \CTMP[15] , \CTMP[14] , \CTMP[13] , \CTMP[12] ,
         \CTMP[11] , \CTMP[10] ;

  HA_0 HA_0 ( .A(A[0]), .B(B[0]), .S(S[0]), .Co(\CTMP[1] ) );
  FA_303 FA_i_2 ( .A(A[1]), .B(B[1]), .Ci(\CTMP[1] ), .S(S[1]), .Co(\CTMP[2] )
         );
  FA_302 FA_i_3 ( .A(A[2]), .B(B[2]), .Ci(\CTMP[2] ), .S(S[2]), .Co(\CTMP[3] )
         );
  FA_301 FA_i_4 ( .A(A[3]), .B(B[3]), .Ci(\CTMP[3] ), .S(S[3]), .Co(\CTMP[4] )
         );
  FA_300 FA_i_5 ( .A(A[4]), .B(B[4]), .Ci(\CTMP[4] ), .S(S[4]), .Co(\CTMP[5] )
         );
  FA_299 FA_i_6 ( .A(A[5]), .B(B[5]), .Ci(\CTMP[5] ), .S(S[5]), .Co(\CTMP[6] )
         );
  FA_298 FA_i_7 ( .A(A[6]), .B(B[6]), .Ci(\CTMP[6] ), .S(S[6]), .Co(\CTMP[7] )
         );
  FA_297 FA_i_8 ( .A(A[7]), .B(B[7]), .Ci(\CTMP[7] ), .S(S[7]), .Co(\CTMP[8] )
         );
  FA_296 FA_i_9 ( .A(A[8]), .B(B[8]), .Ci(\CTMP[8] ), .S(S[8]), .Co(\CTMP[9] )
         );
  FA_295 FA_i_10 ( .A(A[9]), .B(B[9]), .Ci(\CTMP[9] ), .S(S[9]), .Co(
        \CTMP[10] ) );
  FA_294 FA_i_11 ( .A(A[10]), .B(B[10]), .Ci(\CTMP[10] ), .S(S[10]), .Co(
        \CTMP[11] ) );
  FA_293 FA_i_12 ( .A(A[11]), .B(B[11]), .Ci(\CTMP[11] ), .S(S[11]), .Co(
        \CTMP[12] ) );
  FA_292 FA_i_13 ( .A(A[12]), .B(B[12]), .Ci(\CTMP[12] ), .S(S[12]), .Co(
        \CTMP[13] ) );
  FA_291 FA_i_14 ( .A(A[13]), .B(B[13]), .Ci(\CTMP[13] ), .S(S[13]), .Co(
        \CTMP[14] ) );
  FA_290 FA_i_15 ( .A(A[14]), .B(B[14]), .Ci(\CTMP[14] ), .S(S[14]), .Co(
        \CTMP[15] ) );
  FA_289 FA_i_16 ( .A(A[15]), .B(B[15]), .Ci(\CTMP[15] ), .S(S[15]), .Co(
        \CTMP[16] ) );
  FA_288 FA_i_17 ( .A(A[16]), .B(B[16]), .Ci(\CTMP[16] ), .S(S[16]), .Co(
        \CTMP[17] ) );
  FA_287 FA_i_18 ( .A(A[17]), .B(B[17]), .Ci(\CTMP[17] ), .S(S[17]), .Co(
        \CTMP[18] ) );
  FA_286 FA_i_19 ( .A(A[18]), .B(B[18]), .Ci(\CTMP[18] ), .S(S[18]), .Co(
        \CTMP[19] ) );
  FA_285 FA_i_20 ( .A(A[19]), .B(B[19]), .Ci(\CTMP[19] ), .S(S[19]), .Co(Co)
         );
endmodule


module mux5to1_N20 ( A, B, C, D, E, Y, SEL );
  input [19:0] A;
  input [19:0] B;
  input [19:0] C;
  input [19:0] D;
  input [19:0] E;
  output [19:0] Y;
  input [2:0] SEL;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198;

  INV_X1 U1 ( .A(n52), .ZN(n7) );
  BUF_X1 U2 ( .A(n10), .Z(n189) );
  BUF_X1 U3 ( .A(n10), .Z(n188) );
  BUF_X1 U4 ( .A(n11), .Z(n192) );
  BUF_X1 U5 ( .A(n11), .Z(n191) );
  BUF_X1 U6 ( .A(n10), .Z(n190) );
  BUF_X1 U7 ( .A(n11), .Z(n193) );
  INV_X1 U8 ( .A(n50), .ZN(n9) );
  OAI21_X1 U9 ( .B1(SEL[2]), .B2(n51), .A(n52), .ZN(n50) );
  NOR3_X1 U10 ( .A1(n53), .A2(SEL[2]), .A3(n54), .ZN(n10) );
  NOR3_X1 U11 ( .A1(SEL[1]), .A2(SEL[2]), .A3(n54), .ZN(n11) );
  NOR2_X1 U12 ( .A1(SEL[1]), .A2(SEL[0]), .ZN(n51) );
  INV_X1 U13 ( .A(SEL[1]), .ZN(n53) );
  BUF_X1 U14 ( .A(n195), .Z(n197) );
  NOR3_X1 U15 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n53), .ZN(n195) );
  BUF_X1 U16 ( .A(n194), .Z(n196) );
  NOR3_X1 U17 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n53), .ZN(n194) );
  NAND2_X1 U18 ( .A1(SEL[2]), .A2(n51), .ZN(n52) );
  BUF_X1 U19 ( .A(n8), .Z(n198) );
  NOR3_X1 U20 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n53), .ZN(n8) );
  INV_X1 U21 ( .A(SEL[0]), .ZN(n54) );
  NAND2_X1 U22 ( .A1(n28), .A2(n29), .ZN(Y[19]) );
  AOI22_X1 U23 ( .A1(D[19]), .A2(n189), .B1(B[19]), .B2(n192), .ZN(n28) );
  AOI222_X1 U24 ( .A1(E[19]), .A2(n7), .B1(C[19]), .B2(n197), .C1(A[19]), .C2(
        n9), .ZN(n29) );
  NAND2_X1 U25 ( .A1(n30), .A2(n31), .ZN(Y[18]) );
  AOI22_X1 U26 ( .A1(D[18]), .A2(n188), .B1(B[18]), .B2(n191), .ZN(n30) );
  AOI222_X1 U27 ( .A1(E[18]), .A2(n7), .B1(C[18]), .B2(n196), .C1(A[18]), .C2(
        n9), .ZN(n31) );
  NAND2_X1 U28 ( .A1(n32), .A2(n33), .ZN(Y[17]) );
  AOI22_X1 U29 ( .A1(D[17]), .A2(n189), .B1(B[17]), .B2(n192), .ZN(n32) );
  AOI222_X1 U30 ( .A1(E[17]), .A2(n7), .B1(C[17]), .B2(n197), .C1(A[17]), .C2(
        n9), .ZN(n33) );
  NAND2_X1 U31 ( .A1(n34), .A2(n35), .ZN(Y[16]) );
  AOI22_X1 U32 ( .A1(D[16]), .A2(n190), .B1(B[16]), .B2(n193), .ZN(n34) );
  AOI222_X1 U33 ( .A1(E[16]), .A2(n7), .B1(C[16]), .B2(n198), .C1(A[16]), .C2(
        n9), .ZN(n35) );
  NAND2_X1 U34 ( .A1(n36), .A2(n37), .ZN(Y[15]) );
  AOI22_X1 U35 ( .A1(D[15]), .A2(n189), .B1(B[15]), .B2(n192), .ZN(n36) );
  AOI222_X1 U36 ( .A1(E[15]), .A2(n7), .B1(C[15]), .B2(n197), .C1(A[15]), .C2(
        n9), .ZN(n37) );
  NAND2_X1 U37 ( .A1(n38), .A2(n39), .ZN(Y[14]) );
  AOI22_X1 U38 ( .A1(D[14]), .A2(n188), .B1(B[14]), .B2(n191), .ZN(n38) );
  AOI222_X1 U39 ( .A1(E[14]), .A2(n7), .B1(C[14]), .B2(n196), .C1(A[14]), .C2(
        n9), .ZN(n39) );
  NAND2_X1 U40 ( .A1(n40), .A2(n41), .ZN(Y[13]) );
  AOI22_X1 U41 ( .A1(D[13]), .A2(n188), .B1(B[13]), .B2(n191), .ZN(n40) );
  AOI222_X1 U42 ( .A1(E[13]), .A2(n7), .B1(C[13]), .B2(n196), .C1(A[13]), .C2(
        n9), .ZN(n41) );
  NAND2_X1 U43 ( .A1(n42), .A2(n43), .ZN(Y[12]) );
  AOI22_X1 U44 ( .A1(D[12]), .A2(n190), .B1(B[12]), .B2(n193), .ZN(n42) );
  AOI222_X1 U45 ( .A1(E[12]), .A2(n7), .B1(C[12]), .B2(n198), .C1(A[12]), .C2(
        n9), .ZN(n43) );
  NAND2_X1 U46 ( .A1(n44), .A2(n45), .ZN(Y[11]) );
  AOI22_X1 U47 ( .A1(D[11]), .A2(n190), .B1(B[11]), .B2(n193), .ZN(n44) );
  AOI222_X1 U48 ( .A1(E[11]), .A2(n7), .B1(C[11]), .B2(n198), .C1(A[11]), .C2(
        n9), .ZN(n45) );
  NAND2_X1 U49 ( .A1(n46), .A2(n47), .ZN(Y[10]) );
  AOI22_X1 U50 ( .A1(D[10]), .A2(n189), .B1(B[10]), .B2(n192), .ZN(n46) );
  AOI222_X1 U51 ( .A1(E[10]), .A2(n7), .B1(C[10]), .B2(n197), .C1(A[10]), .C2(
        n9), .ZN(n47) );
  NAND2_X1 U52 ( .A1(n5), .A2(n6), .ZN(Y[9]) );
  AOI22_X1 U53 ( .A1(D[9]), .A2(n189), .B1(B[9]), .B2(n192), .ZN(n5) );
  AOI222_X1 U54 ( .A1(E[9]), .A2(n7), .B1(C[9]), .B2(n197), .C1(A[9]), .C2(n9), 
        .ZN(n6) );
  NAND2_X1 U55 ( .A1(n12), .A2(n13), .ZN(Y[8]) );
  AOI22_X1 U56 ( .A1(D[8]), .A2(n188), .B1(B[8]), .B2(n191), .ZN(n12) );
  AOI222_X1 U57 ( .A1(E[8]), .A2(n7), .B1(C[8]), .B2(n196), .C1(A[8]), .C2(n9), 
        .ZN(n13) );
  NAND2_X1 U58 ( .A1(n14), .A2(n15), .ZN(Y[7]) );
  AOI22_X1 U59 ( .A1(D[7]), .A2(n189), .B1(B[7]), .B2(n192), .ZN(n14) );
  AOI222_X1 U60 ( .A1(E[7]), .A2(n7), .B1(C[7]), .B2(n197), .C1(A[7]), .C2(n9), 
        .ZN(n15) );
  NAND2_X1 U61 ( .A1(n16), .A2(n17), .ZN(Y[6]) );
  AOI22_X1 U62 ( .A1(D[6]), .A2(n190), .B1(B[6]), .B2(n193), .ZN(n16) );
  AOI222_X1 U63 ( .A1(E[6]), .A2(n7), .B1(C[6]), .B2(n198), .C1(A[6]), .C2(n9), 
        .ZN(n17) );
  NAND2_X1 U64 ( .A1(n18), .A2(n19), .ZN(Y[5]) );
  AOI22_X1 U65 ( .A1(D[5]), .A2(n189), .B1(B[5]), .B2(n192), .ZN(n18) );
  AOI222_X1 U66 ( .A1(E[5]), .A2(n7), .B1(C[5]), .B2(n197), .C1(A[5]), .C2(n9), 
        .ZN(n19) );
  NAND2_X1 U67 ( .A1(n20), .A2(n21), .ZN(Y[4]) );
  AOI22_X1 U68 ( .A1(D[4]), .A2(n188), .B1(B[4]), .B2(n191), .ZN(n20) );
  AOI222_X1 U69 ( .A1(E[4]), .A2(n7), .B1(C[4]), .B2(n196), .C1(A[4]), .C2(n9), 
        .ZN(n21) );
  NAND2_X1 U70 ( .A1(n22), .A2(n23), .ZN(Y[3]) );
  AOI22_X1 U71 ( .A1(D[3]), .A2(n188), .B1(B[3]), .B2(n191), .ZN(n22) );
  AOI222_X1 U72 ( .A1(E[3]), .A2(n7), .B1(C[3]), .B2(n196), .C1(A[3]), .C2(n9), 
        .ZN(n23) );
  NAND2_X1 U73 ( .A1(n24), .A2(n25), .ZN(Y[2]) );
  AOI22_X1 U74 ( .A1(D[2]), .A2(n190), .B1(B[2]), .B2(n193), .ZN(n24) );
  AOI222_X1 U75 ( .A1(E[2]), .A2(n7), .B1(C[2]), .B2(n198), .C1(A[2]), .C2(n9), 
        .ZN(n25) );
  NAND2_X1 U76 ( .A1(n26), .A2(n27), .ZN(Y[1]) );
  AOI22_X1 U77 ( .A1(D[1]), .A2(n190), .B1(B[1]), .B2(n193), .ZN(n26) );
  AOI222_X1 U78 ( .A1(E[1]), .A2(n7), .B1(C[1]), .B2(n198), .C1(A[1]), .C2(n9), 
        .ZN(n27) );
  NAND2_X1 U79 ( .A1(n48), .A2(n49), .ZN(Y[0]) );
  AOI22_X1 U80 ( .A1(D[0]), .A2(n188), .B1(B[0]), .B2(n191), .ZN(n48) );
  AOI222_X1 U81 ( .A1(E[0]), .A2(n7), .B1(C[0]), .B2(n196), .C1(A[0]), .C2(n9), 
        .ZN(n49) );
endmodule


module mux5to1_N18 ( A, B, C, D, E, Y, SEL );
  input [17:0] A;
  input [17:0] B;
  input [17:0] C;
  input [17:0] D;
  input [17:0] E;
  output [17:0] Y;
  input [2:0] SEL;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47;

  AOI21_X2 U51 ( .B1(n43), .B2(n44), .A(n9), .ZN(n6) );
  XOR2_X1 U63 ( .A(n43), .B(n44), .Z(n24) );
  NOR2_X2 U1 ( .A1(n44), .A2(n43), .ZN(n9) );
  AND3_X1 U2 ( .A1(SEL[0]), .A2(n44), .A3(SEL[1]), .ZN(n7) );
  AND3_X1 U3 ( .A1(n47), .A2(n44), .A3(SEL[0]), .ZN(n5) );
  INV_X1 U4 ( .A(SEL[2]), .ZN(n44) );
  OR2_X1 U5 ( .A1(SEL[0]), .A2(SEL[1]), .ZN(n43) );
  INV_X1 U6 ( .A(SEL[1]), .ZN(n47) );
  NAND2_X1 U7 ( .A1(n27), .A2(n28), .ZN(Y[17]) );
  AOI22_X1 U8 ( .A1(C[17]), .A2(n8), .B1(E[17]), .B2(n9), .ZN(n27) );
  AOI222_X1 U9 ( .A1(B[17]), .A2(n5), .B1(A[17]), .B2(n6), .C1(D[17]), .C2(n7), 
        .ZN(n28) );
  NAND2_X1 U10 ( .A1(n29), .A2(n30), .ZN(Y[16]) );
  AOI22_X1 U11 ( .A1(C[16]), .A2(n8), .B1(E[16]), .B2(n9), .ZN(n29) );
  AOI222_X1 U12 ( .A1(B[16]), .A2(n5), .B1(A[16]), .B2(n6), .C1(D[16]), .C2(n7), .ZN(n30) );
  NAND2_X1 U13 ( .A1(n31), .A2(n32), .ZN(Y[15]) );
  AOI22_X1 U14 ( .A1(C[15]), .A2(n8), .B1(E[15]), .B2(n9), .ZN(n31) );
  AOI222_X1 U15 ( .A1(B[15]), .A2(n5), .B1(A[15]), .B2(n6), .C1(D[15]), .C2(n7), .ZN(n32) );
  NAND2_X1 U16 ( .A1(n33), .A2(n34), .ZN(Y[14]) );
  AOI22_X1 U17 ( .A1(C[14]), .A2(n8), .B1(E[14]), .B2(n9), .ZN(n33) );
  AOI222_X1 U18 ( .A1(B[14]), .A2(n5), .B1(A[14]), .B2(n6), .C1(D[14]), .C2(n7), .ZN(n34) );
  NAND2_X1 U19 ( .A1(n35), .A2(n36), .ZN(Y[13]) );
  AOI22_X1 U20 ( .A1(C[13]), .A2(n8), .B1(E[13]), .B2(n9), .ZN(n35) );
  AOI222_X1 U21 ( .A1(B[13]), .A2(n5), .B1(A[13]), .B2(n6), .C1(D[13]), .C2(n7), .ZN(n36) );
  NAND2_X1 U22 ( .A1(n37), .A2(n38), .ZN(Y[12]) );
  AOI22_X1 U23 ( .A1(C[12]), .A2(n8), .B1(E[12]), .B2(n9), .ZN(n37) );
  AOI222_X1 U24 ( .A1(B[12]), .A2(n5), .B1(A[12]), .B2(n6), .C1(D[12]), .C2(n7), .ZN(n38) );
  NAND2_X1 U25 ( .A1(n39), .A2(n40), .ZN(Y[11]) );
  AOI22_X1 U26 ( .A1(C[11]), .A2(n8), .B1(E[11]), .B2(n9), .ZN(n39) );
  AOI222_X1 U27 ( .A1(B[11]), .A2(n5), .B1(A[11]), .B2(n6), .C1(D[11]), .C2(n7), .ZN(n40) );
  NAND2_X1 U28 ( .A1(n41), .A2(n42), .ZN(Y[10]) );
  AOI22_X1 U29 ( .A1(C[10]), .A2(n8), .B1(E[10]), .B2(n9), .ZN(n41) );
  AOI222_X1 U30 ( .A1(B[10]), .A2(n5), .B1(A[10]), .B2(n6), .C1(D[10]), .C2(n7), .ZN(n42) );
  NAND2_X1 U31 ( .A1(n3), .A2(n4), .ZN(Y[9]) );
  AOI22_X1 U32 ( .A1(C[9]), .A2(n8), .B1(E[9]), .B2(n9), .ZN(n3) );
  AOI222_X1 U33 ( .A1(B[9]), .A2(n5), .B1(A[9]), .B2(n6), .C1(D[9]), .C2(n7), 
        .ZN(n4) );
  NAND2_X1 U34 ( .A1(n10), .A2(n11), .ZN(Y[8]) );
  AOI22_X1 U35 ( .A1(C[8]), .A2(n8), .B1(E[8]), .B2(n9), .ZN(n10) );
  AOI222_X1 U36 ( .A1(B[8]), .A2(n5), .B1(A[8]), .B2(n6), .C1(D[8]), .C2(n7), 
        .ZN(n11) );
  NAND2_X1 U37 ( .A1(n12), .A2(n13), .ZN(Y[7]) );
  AOI22_X1 U38 ( .A1(C[7]), .A2(n8), .B1(E[7]), .B2(n9), .ZN(n12) );
  AOI222_X1 U39 ( .A1(B[7]), .A2(n5), .B1(A[7]), .B2(n6), .C1(D[7]), .C2(n7), 
        .ZN(n13) );
  NAND2_X1 U40 ( .A1(n14), .A2(n15), .ZN(Y[6]) );
  AOI22_X1 U41 ( .A1(C[6]), .A2(n8), .B1(E[6]), .B2(n9), .ZN(n14) );
  AOI222_X1 U42 ( .A1(B[6]), .A2(n5), .B1(A[6]), .B2(n6), .C1(D[6]), .C2(n7), 
        .ZN(n15) );
  NAND2_X1 U43 ( .A1(n16), .A2(n17), .ZN(Y[5]) );
  AOI22_X1 U44 ( .A1(C[5]), .A2(n8), .B1(E[5]), .B2(n9), .ZN(n16) );
  AOI222_X1 U45 ( .A1(B[5]), .A2(n5), .B1(A[5]), .B2(n6), .C1(D[5]), .C2(n7), 
        .ZN(n17) );
  NAND2_X1 U46 ( .A1(n18), .A2(n19), .ZN(Y[4]) );
  AOI22_X1 U47 ( .A1(C[4]), .A2(n8), .B1(E[4]), .B2(n9), .ZN(n18) );
  AOI222_X1 U48 ( .A1(B[4]), .A2(n5), .B1(A[4]), .B2(n6), .C1(D[4]), .C2(n7), 
        .ZN(n19) );
  NAND2_X1 U49 ( .A1(n20), .A2(n21), .ZN(Y[3]) );
  AOI22_X1 U50 ( .A1(C[3]), .A2(n8), .B1(E[3]), .B2(n9), .ZN(n20) );
  AOI222_X1 U52 ( .A1(B[3]), .A2(n5), .B1(A[3]), .B2(n6), .C1(D[3]), .C2(n7), 
        .ZN(n21) );
  NAND2_X1 U53 ( .A1(n25), .A2(n26), .ZN(Y[1]) );
  AOI22_X1 U54 ( .A1(C[1]), .A2(n8), .B1(E[1]), .B2(n9), .ZN(n25) );
  AOI222_X1 U55 ( .A1(B[1]), .A2(n5), .B1(A[1]), .B2(n6), .C1(D[1]), .C2(n7), 
        .ZN(n26) );
  NAND2_X1 U56 ( .A1(n22), .A2(n23), .ZN(Y[2]) );
  AOI22_X1 U57 ( .A1(C[2]), .A2(n8), .B1(E[2]), .B2(n9), .ZN(n22) );
  AOI222_X1 U58 ( .A1(B[2]), .A2(n5), .B1(D[2]), .B2(n7), .C1(A[2]), .C2(n24), 
        .ZN(n23) );
  NAND2_X1 U59 ( .A1(n45), .A2(n46), .ZN(Y[0]) );
  AOI22_X1 U60 ( .A1(C[0]), .A2(n8), .B1(E[0]), .B2(n9), .ZN(n45) );
  AOI222_X1 U61 ( .A1(B[0]), .A2(n5), .B1(D[0]), .B2(n7), .C1(A[0]), .C2(n24), 
        .ZN(n46) );
  NOR3_X4 U62 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n47), .ZN(n8) );
endmodule


module rcas_N16 ( A, B, add_sub, S, Co );
  input [15:0] A;
  input [15:0] B;
  output [15:0] S;
  input add_sub;
  output Co;
  wire   \CTMP[9] , \CTMP[8] , \CTMP[7] , \CTMP[6] , \CTMP[5] , \CTMP[4] ,
         \CTMP[3] , \CTMP[2] , \CTMP[1] , \CTMP[15] , \CTMP[14] , \CTMP[13] ,
         \CTMP[12] , \CTMP[11] , \CTMP[10] ;
  wire   [15:0] Bxor;

  XOR2_X1 U1 ( .A(add_sub), .B(B[9]), .Z(Bxor[9]) );
  XOR2_X1 U2 ( .A(add_sub), .B(B[8]), .Z(Bxor[8]) );
  XOR2_X1 U3 ( .A(add_sub), .B(B[7]), .Z(Bxor[7]) );
  XOR2_X1 U4 ( .A(add_sub), .B(B[6]), .Z(Bxor[6]) );
  XOR2_X1 U5 ( .A(add_sub), .B(B[5]), .Z(Bxor[5]) );
  XOR2_X1 U6 ( .A(add_sub), .B(B[4]), .Z(Bxor[4]) );
  XOR2_X1 U7 ( .A(add_sub), .B(B[3]), .Z(Bxor[3]) );
  XOR2_X1 U8 ( .A(add_sub), .B(B[2]), .Z(Bxor[2]) );
  XOR2_X1 U9 ( .A(add_sub), .B(B[1]), .Z(Bxor[1]) );
  XOR2_X1 U10 ( .A(add_sub), .B(B[15]), .Z(Bxor[15]) );
  XOR2_X1 U11 ( .A(add_sub), .B(B[14]), .Z(Bxor[14]) );
  XOR2_X1 U12 ( .A(add_sub), .B(B[13]), .Z(Bxor[13]) );
  XOR2_X1 U13 ( .A(add_sub), .B(B[12]), .Z(Bxor[12]) );
  XOR2_X1 U14 ( .A(add_sub), .B(B[11]), .Z(Bxor[11]) );
  XOR2_X1 U15 ( .A(add_sub), .B(B[10]), .Z(Bxor[10]) );
  XOR2_X1 U16 ( .A(add_sub), .B(B[0]), .Z(Bxor[0]) );
  FA_0 FA_i_1 ( .A(A[0]), .B(Bxor[0]), .Ci(add_sub), .S(S[0]), .Co(\CTMP[1] )
         );
  FA_318 FA_i_2 ( .A(A[1]), .B(Bxor[1]), .Ci(\CTMP[1] ), .S(S[1]), .Co(
        \CTMP[2] ) );
  FA_317 FA_i_3 ( .A(A[2]), .B(Bxor[2]), .Ci(\CTMP[2] ), .S(S[2]), .Co(
        \CTMP[3] ) );
  FA_316 FA_i_4 ( .A(A[3]), .B(Bxor[3]), .Ci(\CTMP[3] ), .S(S[3]), .Co(
        \CTMP[4] ) );
  FA_315 FA_i_5 ( .A(A[4]), .B(Bxor[4]), .Ci(\CTMP[4] ), .S(S[4]), .Co(
        \CTMP[5] ) );
  FA_314 FA_i_6 ( .A(A[5]), .B(Bxor[5]), .Ci(\CTMP[5] ), .S(S[5]), .Co(
        \CTMP[6] ) );
  FA_313 FA_i_7 ( .A(A[6]), .B(Bxor[6]), .Ci(\CTMP[6] ), .S(S[6]), .Co(
        \CTMP[7] ) );
  FA_312 FA_i_8 ( .A(A[7]), .B(Bxor[7]), .Ci(\CTMP[7] ), .S(S[7]), .Co(
        \CTMP[8] ) );
  FA_311 FA_i_9 ( .A(A[8]), .B(Bxor[8]), .Ci(\CTMP[8] ), .S(S[8]), .Co(
        \CTMP[9] ) );
  FA_310 FA_i_10 ( .A(A[9]), .B(Bxor[9]), .Ci(\CTMP[9] ), .S(S[9]), .Co(
        \CTMP[10] ) );
  FA_309 FA_i_11 ( .A(A[10]), .B(Bxor[10]), .Ci(\CTMP[10] ), .S(S[10]), .Co(
        \CTMP[11] ) );
  FA_308 FA_i_12 ( .A(A[11]), .B(Bxor[11]), .Ci(\CTMP[11] ), .S(S[11]), .Co(
        \CTMP[12] ) );
  FA_307 FA_i_13 ( .A(A[12]), .B(Bxor[12]), .Ci(\CTMP[12] ), .S(S[12]), .Co(
        \CTMP[13] ) );
  FA_306 FA_i_14 ( .A(A[13]), .B(Bxor[13]), .Ci(\CTMP[13] ), .S(S[13]), .Co(
        \CTMP[14] ) );
  FA_305 FA_i_15 ( .A(A[14]), .B(Bxor[14]), .Ci(\CTMP[14] ), .S(S[14]), .Co(
        \CTMP[15] ) );
  FA_304 FA_i_16 ( .A(A[15]), .B(Bxor[15]), .Ci(\CTMP[15] ), .S(S[15]), .Co(Co) );
endmodule


module SHIFTER_GENERIC_N32_DW_rbsh_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \MR_int[1][31] , \MR_int[1][30] , \MR_int[1][29] , \MR_int[1][28] ,
         \MR_int[1][27] , \MR_int[1][26] , \MR_int[1][25] , \MR_int[1][24] ,
         \MR_int[1][23] , \MR_int[1][22] , \MR_int[1][21] , \MR_int[1][20] ,
         \MR_int[1][19] , \MR_int[1][18] , \MR_int[1][17] , \MR_int[1][16] ,
         \MR_int[1][15] , \MR_int[1][14] , \MR_int[1][13] , \MR_int[1][12] ,
         \MR_int[1][11] , \MR_int[1][10] , \MR_int[1][9] , \MR_int[1][8] ,
         \MR_int[1][7] , \MR_int[1][6] , \MR_int[1][5] , \MR_int[1][4] ,
         \MR_int[1][3] , \MR_int[1][2] , \MR_int[1][1] , \MR_int[1][0] ,
         \MR_int[2][31] , \MR_int[2][30] , \MR_int[2][29] , \MR_int[2][28] ,
         \MR_int[2][27] , \MR_int[2][26] , \MR_int[2][25] , \MR_int[2][24] ,
         \MR_int[2][23] , \MR_int[2][22] , \MR_int[2][21] , \MR_int[2][20] ,
         \MR_int[2][19] , \MR_int[2][18] , \MR_int[2][17] , \MR_int[2][16] ,
         \MR_int[2][15] , \MR_int[2][14] , \MR_int[2][13] , \MR_int[2][12] ,
         \MR_int[2][11] , \MR_int[2][10] , \MR_int[2][9] , \MR_int[2][8] ,
         \MR_int[2][7] , \MR_int[2][6] , \MR_int[2][5] , \MR_int[2][4] ,
         \MR_int[2][3] , \MR_int[2][2] , \MR_int[2][1] , \MR_int[2][0] ,
         \MR_int[3][31] , \MR_int[3][30] , \MR_int[3][29] , \MR_int[3][28] ,
         \MR_int[3][27] , \MR_int[3][26] , \MR_int[3][25] , \MR_int[3][24] ,
         \MR_int[3][23] , \MR_int[3][22] , \MR_int[3][21] , \MR_int[3][20] ,
         \MR_int[3][19] , \MR_int[3][18] , \MR_int[3][17] , \MR_int[3][16] ,
         \MR_int[3][15] , \MR_int[3][14] , \MR_int[3][13] , \MR_int[3][12] ,
         \MR_int[3][11] , \MR_int[3][10] , \MR_int[3][9] , \MR_int[3][8] ,
         \MR_int[3][7] , \MR_int[3][6] , \MR_int[3][5] , \MR_int[3][4] ,
         \MR_int[3][3] , \MR_int[3][2] , \MR_int[3][1] , \MR_int[3][0] ,
         \MR_int[4][31] , \MR_int[4][30] , \MR_int[4][29] , \MR_int[4][28] ,
         \MR_int[4][27] , \MR_int[4][26] , \MR_int[4][25] , \MR_int[4][24] ,
         \MR_int[4][23] , \MR_int[4][22] , \MR_int[4][21] , \MR_int[4][20] ,
         \MR_int[4][19] , \MR_int[4][18] , \MR_int[4][17] , \MR_int[4][16] ,
         \MR_int[4][15] , \MR_int[4][14] , \MR_int[4][13] , \MR_int[4][12] ,
         \MR_int[4][11] , \MR_int[4][10] , \MR_int[4][9] , \MR_int[4][8] ,
         \MR_int[4][7] , \MR_int[4][6] , \MR_int[4][5] , \MR_int[4][4] ,
         \MR_int[4][3] , \MR_int[4][2] , \MR_int[4][1] , \MR_int[4][0] , n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138;

  MUX2_X1 M1_4_31 ( .A(\MR_int[4][31] ), .B(\MR_int[4][15] ), .S(n137), .Z(
        B[31]) );
  MUX2_X1 M1_4_30 ( .A(\MR_int[4][30] ), .B(\MR_int[4][14] ), .S(n137), .Z(
        B[30]) );
  MUX2_X1 M1_4_29 ( .A(\MR_int[4][29] ), .B(\MR_int[4][13] ), .S(n137), .Z(
        B[29]) );
  MUX2_X1 M1_4_28 ( .A(\MR_int[4][28] ), .B(\MR_int[4][12] ), .S(n137), .Z(
        B[28]) );
  MUX2_X1 M1_4_27 ( .A(\MR_int[4][27] ), .B(\MR_int[4][11] ), .S(n137), .Z(
        B[27]) );
  MUX2_X1 M1_4_26 ( .A(\MR_int[4][26] ), .B(\MR_int[4][10] ), .S(n137), .Z(
        B[26]) );
  MUX2_X1 M1_4_25 ( .A(\MR_int[4][25] ), .B(\MR_int[4][9] ), .S(n137), .Z(
        B[25]) );
  MUX2_X1 M1_4_24 ( .A(\MR_int[4][24] ), .B(\MR_int[4][8] ), .S(n137), .Z(
        B[24]) );
  MUX2_X1 M1_4_23 ( .A(\MR_int[4][23] ), .B(\MR_int[4][7] ), .S(n137), .Z(
        B[23]) );
  MUX2_X1 M1_4_22 ( .A(\MR_int[4][22] ), .B(\MR_int[4][6] ), .S(n136), .Z(
        B[22]) );
  MUX2_X1 M1_4_21 ( .A(\MR_int[4][21] ), .B(\MR_int[4][5] ), .S(n136), .Z(
        B[21]) );
  MUX2_X1 M1_4_20 ( .A(\MR_int[4][20] ), .B(\MR_int[4][4] ), .S(n136), .Z(
        B[20]) );
  MUX2_X1 M1_4_19 ( .A(\MR_int[4][19] ), .B(\MR_int[4][3] ), .S(n136), .Z(
        B[19]) );
  MUX2_X1 M1_4_18 ( .A(\MR_int[4][18] ), .B(\MR_int[4][2] ), .S(n136), .Z(
        B[18]) );
  MUX2_X1 M1_4_17 ( .A(\MR_int[4][17] ), .B(\MR_int[4][1] ), .S(n136), .Z(
        B[17]) );
  MUX2_X1 M1_4_16 ( .A(\MR_int[4][16] ), .B(\MR_int[4][0] ), .S(n136), .Z(
        B[16]) );
  MUX2_X1 M1_4_15 ( .A(\MR_int[4][15] ), .B(\MR_int[4][31] ), .S(n136), .Z(
        B[15]) );
  MUX2_X1 M1_4_14 ( .A(\MR_int[4][14] ), .B(\MR_int[4][30] ), .S(n136), .Z(
        B[14]) );
  MUX2_X1 M1_4_13 ( .A(\MR_int[4][13] ), .B(\MR_int[4][29] ), .S(n136), .Z(
        B[13]) );
  MUX2_X1 M1_4_12 ( .A(\MR_int[4][12] ), .B(\MR_int[4][28] ), .S(n136), .Z(
        B[12]) );
  MUX2_X1 M1_4_11 ( .A(\MR_int[4][11] ), .B(\MR_int[4][27] ), .S(n136), .Z(
        B[11]) );
  MUX2_X1 M1_4_10 ( .A(\MR_int[4][10] ), .B(\MR_int[4][26] ), .S(n138), .Z(
        B[10]) );
  MUX2_X1 M1_4_9 ( .A(\MR_int[4][9] ), .B(\MR_int[4][25] ), .S(n137), .Z(B[9])
         );
  MUX2_X1 M1_4_8 ( .A(\MR_int[4][8] ), .B(\MR_int[4][24] ), .S(n138), .Z(B[8])
         );
  MUX2_X1 M1_4_7 ( .A(\MR_int[4][7] ), .B(\MR_int[4][23] ), .S(n138), .Z(B[7])
         );
  MUX2_X1 M1_4_6 ( .A(\MR_int[4][6] ), .B(\MR_int[4][22] ), .S(n138), .Z(B[6])
         );
  MUX2_X1 M1_4_5 ( .A(\MR_int[4][5] ), .B(\MR_int[4][21] ), .S(n137), .Z(B[5])
         );
  MUX2_X1 M1_4_4 ( .A(\MR_int[4][4] ), .B(\MR_int[4][20] ), .S(n138), .Z(B[4])
         );
  MUX2_X1 M1_4_3 ( .A(\MR_int[4][3] ), .B(\MR_int[4][19] ), .S(n138), .Z(B[3])
         );
  MUX2_X1 M1_4_2 ( .A(\MR_int[4][2] ), .B(\MR_int[4][18] ), .S(n138), .Z(B[2])
         );
  MUX2_X1 M1_4_1 ( .A(\MR_int[4][1] ), .B(\MR_int[4][17] ), .S(n138), .Z(B[1])
         );
  MUX2_X1 M1_4_0 ( .A(\MR_int[4][0] ), .B(\MR_int[4][16] ), .S(n137), .Z(B[0])
         );
  MUX2_X1 M1_3_31_0 ( .A(\MR_int[3][31] ), .B(\MR_int[3][7] ), .S(n134), .Z(
        \MR_int[4][31] ) );
  MUX2_X1 M1_3_30_0 ( .A(\MR_int[3][30] ), .B(\MR_int[3][6] ), .S(n134), .Z(
        \MR_int[4][30] ) );
  MUX2_X1 M1_3_29_0 ( .A(\MR_int[3][29] ), .B(\MR_int[3][5] ), .S(n134), .Z(
        \MR_int[4][29] ) );
  MUX2_X1 M1_3_28_0 ( .A(\MR_int[3][28] ), .B(\MR_int[3][4] ), .S(n134), .Z(
        \MR_int[4][28] ) );
  MUX2_X1 M1_3_27_0 ( .A(\MR_int[3][27] ), .B(\MR_int[3][3] ), .S(n134), .Z(
        \MR_int[4][27] ) );
  MUX2_X1 M1_3_26_0 ( .A(\MR_int[3][26] ), .B(\MR_int[3][2] ), .S(n134), .Z(
        \MR_int[4][26] ) );
  MUX2_X1 M1_3_25_0 ( .A(\MR_int[3][25] ), .B(\MR_int[3][1] ), .S(n134), .Z(
        \MR_int[4][25] ) );
  MUX2_X1 M1_3_24_0 ( .A(\MR_int[3][24] ), .B(\MR_int[3][0] ), .S(n133), .Z(
        \MR_int[4][24] ) );
  MUX2_X1 M1_3_23_0 ( .A(\MR_int[3][23] ), .B(\MR_int[3][31] ), .S(n133), .Z(
        \MR_int[4][23] ) );
  MUX2_X1 M1_3_22_0 ( .A(\MR_int[3][22] ), .B(\MR_int[3][30] ), .S(n133), .Z(
        \MR_int[4][22] ) );
  MUX2_X1 M1_3_21_0 ( .A(\MR_int[3][21] ), .B(\MR_int[3][29] ), .S(n133), .Z(
        \MR_int[4][21] ) );
  MUX2_X1 M1_3_20_0 ( .A(\MR_int[3][20] ), .B(\MR_int[3][28] ), .S(n133), .Z(
        \MR_int[4][20] ) );
  MUX2_X1 M1_3_19_0 ( .A(\MR_int[3][19] ), .B(\MR_int[3][27] ), .S(n133), .Z(
        \MR_int[4][19] ) );
  MUX2_X1 M1_3_18_0 ( .A(\MR_int[3][18] ), .B(\MR_int[3][26] ), .S(n133), .Z(
        \MR_int[4][18] ) );
  MUX2_X1 M1_3_17_0 ( .A(\MR_int[3][17] ), .B(\MR_int[3][25] ), .S(n135), .Z(
        \MR_int[4][17] ) );
  MUX2_X1 M1_3_16_0 ( .A(\MR_int[3][16] ), .B(\MR_int[3][24] ), .S(n135), .Z(
        \MR_int[4][16] ) );
  MUX2_X1 M1_3_15_0 ( .A(\MR_int[3][15] ), .B(\MR_int[3][23] ), .S(n135), .Z(
        \MR_int[4][15] ) );
  MUX2_X1 M1_3_14_0 ( .A(\MR_int[3][14] ), .B(\MR_int[3][22] ), .S(n134), .Z(
        \MR_int[4][14] ) );
  MUX2_X1 M1_3_13_0 ( .A(\MR_int[3][13] ), .B(\MR_int[3][21] ), .S(n134), .Z(
        \MR_int[4][13] ) );
  MUX2_X1 M1_3_12_0 ( .A(\MR_int[3][12] ), .B(\MR_int[3][20] ), .S(n134), .Z(
        \MR_int[4][12] ) );
  MUX2_X1 M1_3_11_0 ( .A(\MR_int[3][11] ), .B(\MR_int[3][19] ), .S(n134), .Z(
        \MR_int[4][11] ) );
  MUX2_X1 M1_3_10_0 ( .A(\MR_int[3][10] ), .B(\MR_int[3][18] ), .S(n133), .Z(
        \MR_int[4][10] ) );
  MUX2_X1 M1_3_9_0 ( .A(\MR_int[3][9] ), .B(\MR_int[3][17] ), .S(n133), .Z(
        \MR_int[4][9] ) );
  MUX2_X1 M1_3_8_0 ( .A(\MR_int[3][8] ), .B(\MR_int[3][16] ), .S(n135), .Z(
        \MR_int[4][8] ) );
  MUX2_X1 M1_3_7 ( .A(\MR_int[3][7] ), .B(\MR_int[3][15] ), .S(n133), .Z(
        \MR_int[4][7] ) );
  MUX2_X1 M1_3_6 ( .A(\MR_int[3][6] ), .B(\MR_int[3][14] ), .S(n133), .Z(
        \MR_int[4][6] ) );
  MUX2_X1 M1_3_5 ( .A(\MR_int[3][5] ), .B(\MR_int[3][13] ), .S(n134), .Z(
        \MR_int[4][5] ) );
  MUX2_X1 M1_3_4 ( .A(\MR_int[3][4] ), .B(\MR_int[3][12] ), .S(n133), .Z(
        \MR_int[4][4] ) );
  MUX2_X1 M1_3_3 ( .A(\MR_int[3][3] ), .B(\MR_int[3][11] ), .S(n135), .Z(
        \MR_int[4][3] ) );
  MUX2_X1 M1_3_2 ( .A(\MR_int[3][2] ), .B(\MR_int[3][10] ), .S(n135), .Z(
        \MR_int[4][2] ) );
  MUX2_X1 M1_3_1 ( .A(\MR_int[3][1] ), .B(\MR_int[3][9] ), .S(n135), .Z(
        \MR_int[4][1] ) );
  MUX2_X1 M1_3_0 ( .A(\MR_int[3][0] ), .B(\MR_int[3][8] ), .S(n135), .Z(
        \MR_int[4][0] ) );
  MUX2_X1 M1_2_31_0 ( .A(\MR_int[2][31] ), .B(\MR_int[2][3] ), .S(n132), .Z(
        \MR_int[3][31] ) );
  MUX2_X1 M1_2_30_0 ( .A(\MR_int[2][30] ), .B(\MR_int[2][2] ), .S(n132), .Z(
        \MR_int[3][30] ) );
  MUX2_X1 M1_2_29_0 ( .A(\MR_int[2][29] ), .B(\MR_int[2][1] ), .S(n132), .Z(
        \MR_int[3][29] ) );
  MUX2_X1 M1_2_28_0 ( .A(\MR_int[2][28] ), .B(\MR_int[2][0] ), .S(n132), .Z(
        \MR_int[3][28] ) );
  MUX2_X1 M1_2_27_0 ( .A(\MR_int[2][27] ), .B(\MR_int[2][31] ), .S(n132), .Z(
        \MR_int[3][27] ) );
  MUX2_X1 M1_2_26_0 ( .A(\MR_int[2][26] ), .B(\MR_int[2][30] ), .S(n132), .Z(
        \MR_int[3][26] ) );
  MUX2_X1 M1_2_25_0 ( .A(\MR_int[2][25] ), .B(\MR_int[2][29] ), .S(n132), .Z(
        \MR_int[3][25] ) );
  MUX2_X1 M1_2_24_0 ( .A(\MR_int[2][24] ), .B(\MR_int[2][28] ), .S(n130), .Z(
        \MR_int[3][24] ) );
  MUX2_X1 M1_2_23_0 ( .A(\MR_int[2][23] ), .B(\MR_int[2][27] ), .S(n130), .Z(
        \MR_int[3][23] ) );
  MUX2_X1 M1_2_22_0 ( .A(\MR_int[2][22] ), .B(\MR_int[2][26] ), .S(n130), .Z(
        \MR_int[3][22] ) );
  MUX2_X1 M1_2_21_0 ( .A(\MR_int[2][21] ), .B(\MR_int[2][25] ), .S(n130), .Z(
        \MR_int[3][21] ) );
  MUX2_X1 M1_2_20_0 ( .A(\MR_int[2][20] ), .B(\MR_int[2][24] ), .S(n130), .Z(
        \MR_int[3][20] ) );
  MUX2_X1 M1_2_19_0 ( .A(\MR_int[2][19] ), .B(\MR_int[2][23] ), .S(n130), .Z(
        \MR_int[3][19] ) );
  MUX2_X1 M1_2_18_0 ( .A(\MR_int[2][18] ), .B(\MR_int[2][22] ), .S(n131), .Z(
        \MR_int[3][18] ) );
  MUX2_X1 M1_2_17_0 ( .A(\MR_int[2][17] ), .B(\MR_int[2][21] ), .S(n132), .Z(
        \MR_int[3][17] ) );
  MUX2_X1 M1_2_16_0 ( .A(\MR_int[2][16] ), .B(\MR_int[2][20] ), .S(n130), .Z(
        \MR_int[3][16] ) );
  MUX2_X1 M1_2_15_0 ( .A(\MR_int[2][15] ), .B(\MR_int[2][19] ), .S(n130), .Z(
        \MR_int[3][15] ) );
  MUX2_X1 M1_2_14_0 ( .A(\MR_int[2][14] ), .B(\MR_int[2][18] ), .S(n130), .Z(
        \MR_int[3][14] ) );
  MUX2_X1 M1_2_13_0 ( .A(\MR_int[2][13] ), .B(\MR_int[2][17] ), .S(n130), .Z(
        \MR_int[3][13] ) );
  MUX2_X1 M1_2_12_0 ( .A(\MR_int[2][12] ), .B(\MR_int[2][16] ), .S(n130), .Z(
        \MR_int[3][12] ) );
  MUX2_X1 M1_2_11_0 ( .A(\MR_int[2][11] ), .B(\MR_int[2][15] ), .S(n130), .Z(
        \MR_int[3][11] ) );
  MUX2_X1 M1_2_10_0 ( .A(\MR_int[2][10] ), .B(\MR_int[2][14] ), .S(n131), .Z(
        \MR_int[3][10] ) );
  MUX2_X1 M1_2_9_0 ( .A(\MR_int[2][9] ), .B(\MR_int[2][13] ), .S(n131), .Z(
        \MR_int[3][9] ) );
  MUX2_X1 M1_2_8_0 ( .A(\MR_int[2][8] ), .B(\MR_int[2][12] ), .S(n131), .Z(
        \MR_int[3][8] ) );
  MUX2_X1 M1_2_7_0 ( .A(\MR_int[2][7] ), .B(\MR_int[2][11] ), .S(n131), .Z(
        \MR_int[3][7] ) );
  MUX2_X1 M1_2_6_0 ( .A(\MR_int[2][6] ), .B(\MR_int[2][10] ), .S(n131), .Z(
        \MR_int[3][6] ) );
  MUX2_X1 M1_2_5_0 ( .A(\MR_int[2][5] ), .B(\MR_int[2][9] ), .S(n131), .Z(
        \MR_int[3][5] ) );
  MUX2_X1 M1_2_4_0 ( .A(\MR_int[2][4] ), .B(\MR_int[2][8] ), .S(n131), .Z(
        \MR_int[3][4] ) );
  MUX2_X1 M1_2_3 ( .A(\MR_int[2][3] ), .B(\MR_int[2][7] ), .S(n131), .Z(
        \MR_int[3][3] ) );
  MUX2_X1 M1_2_2 ( .A(\MR_int[2][2] ), .B(\MR_int[2][6] ), .S(n131), .Z(
        \MR_int[3][2] ) );
  MUX2_X1 M1_2_1 ( .A(\MR_int[2][1] ), .B(\MR_int[2][5] ), .S(n131), .Z(
        \MR_int[3][1] ) );
  MUX2_X1 M1_2_0 ( .A(\MR_int[2][0] ), .B(\MR_int[2][4] ), .S(n131), .Z(
        \MR_int[3][0] ) );
  MUX2_X1 M1_1_31_0 ( .A(\MR_int[1][31] ), .B(\MR_int[1][1] ), .S(n128), .Z(
        \MR_int[2][31] ) );
  MUX2_X1 M1_1_30_0 ( .A(\MR_int[1][30] ), .B(\MR_int[1][0] ), .S(n128), .Z(
        \MR_int[2][30] ) );
  MUX2_X1 M1_1_29_0 ( .A(\MR_int[1][29] ), .B(\MR_int[1][31] ), .S(n128), .Z(
        \MR_int[2][29] ) );
  MUX2_X1 M1_1_28_0 ( .A(\MR_int[1][28] ), .B(\MR_int[1][30] ), .S(n128), .Z(
        \MR_int[2][28] ) );
  MUX2_X1 M1_1_27_0 ( .A(\MR_int[1][27] ), .B(\MR_int[1][29] ), .S(n128), .Z(
        \MR_int[2][27] ) );
  MUX2_X1 M1_1_26_0 ( .A(\MR_int[1][26] ), .B(\MR_int[1][28] ), .S(n128), .Z(
        \MR_int[2][26] ) );
  MUX2_X1 M1_1_25_0 ( .A(\MR_int[1][25] ), .B(\MR_int[1][27] ), .S(n128), .Z(
        \MR_int[2][25] ) );
  MUX2_X1 M1_1_24_0 ( .A(\MR_int[1][24] ), .B(\MR_int[1][26] ), .S(n129), .Z(
        \MR_int[2][24] ) );
  MUX2_X1 M1_1_23_0 ( .A(\MR_int[1][23] ), .B(\MR_int[1][25] ), .S(n128), .Z(
        \MR_int[2][23] ) );
  MUX2_X1 M1_1_22_0 ( .A(\MR_int[1][22] ), .B(\MR_int[1][24] ), .S(n128), .Z(
        \MR_int[2][22] ) );
  MUX2_X1 M1_1_21_0 ( .A(\MR_int[1][21] ), .B(\MR_int[1][23] ), .S(n128), .Z(
        \MR_int[2][21] ) );
  MUX2_X1 M1_1_20_0 ( .A(\MR_int[1][20] ), .B(\MR_int[1][22] ), .S(n127), .Z(
        \MR_int[2][20] ) );
  MUX2_X1 M1_1_19_0 ( .A(\MR_int[1][19] ), .B(\MR_int[1][21] ), .S(n128), .Z(
        \MR_int[2][19] ) );
  MUX2_X1 M1_1_18_0 ( .A(\MR_int[1][18] ), .B(\MR_int[1][20] ), .S(n127), .Z(
        \MR_int[2][18] ) );
  MUX2_X1 M1_1_17_0 ( .A(\MR_int[1][17] ), .B(\MR_int[1][19] ), .S(n127), .Z(
        \MR_int[2][17] ) );
  MUX2_X1 M1_1_16_0 ( .A(\MR_int[1][16] ), .B(\MR_int[1][18] ), .S(n127), .Z(
        \MR_int[2][16] ) );
  MUX2_X1 M1_1_15_0 ( .A(\MR_int[1][15] ), .B(\MR_int[1][17] ), .S(n127), .Z(
        \MR_int[2][15] ) );
  MUX2_X1 M1_1_14_0 ( .A(\MR_int[1][14] ), .B(\MR_int[1][16] ), .S(n127), .Z(
        \MR_int[2][14] ) );
  MUX2_X1 M1_1_13_0 ( .A(\MR_int[1][13] ), .B(\MR_int[1][15] ), .S(n127), .Z(
        \MR_int[2][13] ) );
  MUX2_X1 M1_1_12_0 ( .A(\MR_int[1][12] ), .B(\MR_int[1][14] ), .S(n127), .Z(
        \MR_int[2][12] ) );
  MUX2_X1 M1_1_11_0 ( .A(\MR_int[1][11] ), .B(\MR_int[1][13] ), .S(n127), .Z(
        \MR_int[2][11] ) );
  MUX2_X1 M1_1_10_0 ( .A(\MR_int[1][10] ), .B(\MR_int[1][12] ), .S(n129), .Z(
        \MR_int[2][10] ) );
  MUX2_X1 M1_1_9_0 ( .A(\MR_int[1][9] ), .B(\MR_int[1][11] ), .S(n129), .Z(
        \MR_int[2][9] ) );
  MUX2_X1 M1_1_8_0 ( .A(\MR_int[1][8] ), .B(\MR_int[1][10] ), .S(n129), .Z(
        \MR_int[2][8] ) );
  MUX2_X1 M1_1_7_0 ( .A(\MR_int[1][7] ), .B(\MR_int[1][9] ), .S(n129), .Z(
        \MR_int[2][7] ) );
  MUX2_X1 M1_1_6_0 ( .A(\MR_int[1][6] ), .B(\MR_int[1][8] ), .S(n129), .Z(
        \MR_int[2][6] ) );
  MUX2_X1 M1_1_5_0 ( .A(\MR_int[1][5] ), .B(\MR_int[1][7] ), .S(n129), .Z(
        \MR_int[2][5] ) );
  MUX2_X1 M1_1_4_0 ( .A(\MR_int[1][4] ), .B(\MR_int[1][6] ), .S(n129), .Z(
        \MR_int[2][4] ) );
  MUX2_X1 M1_1_3_0 ( .A(\MR_int[1][3] ), .B(\MR_int[1][5] ), .S(n128), .Z(
        \MR_int[2][3] ) );
  MUX2_X1 M1_1_2_0 ( .A(\MR_int[1][2] ), .B(\MR_int[1][4] ), .S(n127), .Z(
        \MR_int[2][2] ) );
  MUX2_X1 M1_1_1 ( .A(\MR_int[1][1] ), .B(\MR_int[1][3] ), .S(n127), .Z(
        \MR_int[2][1] ) );
  MUX2_X1 M1_1_0 ( .A(\MR_int[1][0] ), .B(\MR_int[1][2] ), .S(n127), .Z(
        \MR_int[2][0] ) );
  MUX2_X1 M1_0_31_0 ( .A(A[31]), .B(A[0]), .S(n125), .Z(\MR_int[1][31] ) );
  MUX2_X1 M1_0_30_0 ( .A(A[30]), .B(A[31]), .S(n125), .Z(\MR_int[1][30] ) );
  MUX2_X1 M1_0_29_0 ( .A(A[29]), .B(A[30]), .S(n125), .Z(\MR_int[1][29] ) );
  MUX2_X1 M1_0_28_0 ( .A(A[28]), .B(A[29]), .S(n125), .Z(\MR_int[1][28] ) );
  MUX2_X1 M1_0_27_0 ( .A(A[27]), .B(A[28]), .S(n125), .Z(\MR_int[1][27] ) );
  MUX2_X1 M1_0_26_0 ( .A(A[26]), .B(A[27]), .S(n125), .Z(\MR_int[1][26] ) );
  MUX2_X1 M1_0_25_0 ( .A(A[25]), .B(A[26]), .S(n125), .Z(\MR_int[1][25] ) );
  MUX2_X1 M1_0_24_0 ( .A(A[24]), .B(A[25]), .S(n125), .Z(\MR_int[1][24] ) );
  MUX2_X1 M1_0_23_0 ( .A(A[23]), .B(A[24]), .S(n124), .Z(\MR_int[1][23] ) );
  MUX2_X1 M1_0_22_0 ( .A(A[22]), .B(A[23]), .S(n124), .Z(\MR_int[1][22] ) );
  MUX2_X1 M1_0_21_0 ( .A(A[21]), .B(A[22]), .S(n124), .Z(\MR_int[1][21] ) );
  MUX2_X1 M1_0_20_0 ( .A(A[20]), .B(A[21]), .S(n124), .Z(\MR_int[1][20] ) );
  MUX2_X1 M1_0_19_0 ( .A(A[19]), .B(A[20]), .S(n125), .Z(\MR_int[1][19] ) );
  MUX2_X1 M1_0_18_0 ( .A(A[18]), .B(A[19]), .S(n124), .Z(\MR_int[1][18] ) );
  MUX2_X1 M1_0_17_0 ( .A(A[17]), .B(A[18]), .S(n124), .Z(\MR_int[1][17] ) );
  MUX2_X1 M1_0_16_0 ( .A(A[16]), .B(A[17]), .S(n124), .Z(\MR_int[1][16] ) );
  MUX2_X1 M1_0_15_0 ( .A(A[15]), .B(A[16]), .S(n124), .Z(\MR_int[1][15] ) );
  MUX2_X1 M1_0_14_0 ( .A(A[14]), .B(A[15]), .S(n124), .Z(\MR_int[1][14] ) );
  MUX2_X1 M1_0_13_0 ( .A(A[13]), .B(A[14]), .S(n124), .Z(\MR_int[1][13] ) );
  MUX2_X1 M1_0_12_0 ( .A(A[12]), .B(A[13]), .S(n124), .Z(\MR_int[1][12] ) );
  MUX2_X1 M1_0_11_0 ( .A(A[11]), .B(A[12]), .S(n124), .Z(\MR_int[1][11] ) );
  MUX2_X1 M1_0_10_0 ( .A(A[10]), .B(A[11]), .S(n126), .Z(\MR_int[1][10] ) );
  MUX2_X1 M1_0_9_0 ( .A(A[9]), .B(A[10]), .S(n126), .Z(\MR_int[1][9] ) );
  MUX2_X1 M1_0_8_0 ( .A(A[8]), .B(A[9]), .S(n126), .Z(\MR_int[1][8] ) );
  MUX2_X1 M1_0_7_0 ( .A(A[7]), .B(A[8]), .S(n126), .Z(\MR_int[1][7] ) );
  MUX2_X1 M1_0_6_0 ( .A(A[6]), .B(A[7]), .S(n126), .Z(\MR_int[1][6] ) );
  MUX2_X1 M1_0_5_0 ( .A(A[5]), .B(A[6]), .S(n126), .Z(\MR_int[1][5] ) );
  MUX2_X1 M1_0_4_0 ( .A(A[4]), .B(A[5]), .S(n125), .Z(\MR_int[1][4] ) );
  MUX2_X1 M1_0_3_0 ( .A(A[3]), .B(A[4]), .S(n126), .Z(\MR_int[1][3] ) );
  MUX2_X1 M1_0_2_0 ( .A(A[2]), .B(A[3]), .S(n126), .Z(\MR_int[1][2] ) );
  MUX2_X1 M1_0_1_0 ( .A(A[1]), .B(A[2]), .S(n125), .Z(\MR_int[1][1] ) );
  MUX2_X1 M1_0_0 ( .A(A[0]), .B(A[1]), .S(n125), .Z(\MR_int[1][0] ) );
  BUF_X1 U2 ( .A(SH[1]), .Z(n127) );
  BUF_X1 U3 ( .A(SH[1]), .Z(n128) );
  BUF_X1 U4 ( .A(SH[3]), .Z(n133) );
  BUF_X1 U5 ( .A(SH[3]), .Z(n134) );
  BUF_X1 U6 ( .A(SH[4]), .Z(n136) );
  BUF_X1 U7 ( .A(SH[4]), .Z(n137) );
  BUF_X1 U8 ( .A(SH[1]), .Z(n129) );
  BUF_X1 U9 ( .A(SH[3]), .Z(n135) );
  BUF_X1 U10 ( .A(SH[4]), .Z(n138) );
  BUF_X1 U11 ( .A(SH[0]), .Z(n124) );
  BUF_X1 U12 ( .A(SH[0]), .Z(n125) );
  BUF_X1 U13 ( .A(SH[2]), .Z(n130) );
  BUF_X1 U14 ( .A(SH[2]), .Z(n131) );
  BUF_X1 U15 ( .A(SH[0]), .Z(n126) );
  BUF_X1 U16 ( .A(SH[2]), .Z(n132) );
endmodule


module SHIFTER_GENERIC_N32_DW_lbsh_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] , \ML_int[1][28] ,
         \ML_int[1][27] , \ML_int[1][26] , \ML_int[1][25] , \ML_int[1][24] ,
         \ML_int[1][23] , \ML_int[1][22] , \ML_int[1][21] , \ML_int[1][20] ,
         \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][31] , \ML_int[2][30] , \ML_int[2][29] , \ML_int[2][28] ,
         \ML_int[2][27] , \ML_int[2][26] , \ML_int[2][25] , \ML_int[2][24] ,
         \ML_int[2][23] , \ML_int[2][22] , \ML_int[2][21] , \ML_int[2][20] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][31] , \ML_int[3][30] , \ML_int[3][29] , \ML_int[3][28] ,
         \ML_int[3][27] , \ML_int[3][26] , \ML_int[3][25] , \ML_int[3][24] ,
         \ML_int[3][23] , \ML_int[3][22] , \ML_int[3][21] , \ML_int[3][20] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[3][3] , \ML_int[3][2] , \ML_int[3][1] , \ML_int[3][0] ,
         \ML_int[4][31] , \ML_int[4][30] , \ML_int[4][29] , \ML_int[4][28] ,
         \ML_int[4][27] , \ML_int[4][26] , \ML_int[4][25] , \ML_int[4][24] ,
         \ML_int[4][23] , \ML_int[4][22] , \ML_int[4][21] , \ML_int[4][20] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][16] ,
         \ML_int[4][15] , \ML_int[4][14] , \ML_int[4][13] , \ML_int[4][12] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[4][7] , \ML_int[4][6] , \ML_int[4][5] , \ML_int[4][4] ,
         \ML_int[4][3] , \ML_int[4][2] , \ML_int[4][1] , \ML_int[4][0] , n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139;

  MUX2_X1 M1_4_31 ( .A(\ML_int[4][31] ), .B(\ML_int[4][15] ), .S(n138), .Z(
        B[31]) );
  MUX2_X1 M1_4_30 ( .A(\ML_int[4][30] ), .B(\ML_int[4][14] ), .S(n138), .Z(
        B[30]) );
  MUX2_X1 M1_4_29 ( .A(\ML_int[4][29] ), .B(\ML_int[4][13] ), .S(n138), .Z(
        B[29]) );
  MUX2_X1 M1_4_28 ( .A(\ML_int[4][28] ), .B(\ML_int[4][12] ), .S(n138), .Z(
        B[28]) );
  MUX2_X1 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S(n138), .Z(
        B[27]) );
  MUX2_X1 M1_4_26 ( .A(\ML_int[4][26] ), .B(\ML_int[4][10] ), .S(n138), .Z(
        B[26]) );
  MUX2_X1 M1_4_25 ( .A(\ML_int[4][25] ), .B(\ML_int[4][9] ), .S(n138), .Z(
        B[25]) );
  MUX2_X1 M1_4_24 ( .A(\ML_int[4][24] ), .B(\ML_int[4][8] ), .S(n138), .Z(
        B[24]) );
  MUX2_X1 M1_4_23 ( .A(\ML_int[4][23] ), .B(\ML_int[4][7] ), .S(n138), .Z(
        B[23]) );
  MUX2_X1 M1_4_22 ( .A(\ML_int[4][22] ), .B(\ML_int[4][6] ), .S(n138), .Z(
        B[22]) );
  MUX2_X1 M1_4_21 ( .A(\ML_int[4][21] ), .B(\ML_int[4][5] ), .S(n138), .Z(
        B[21]) );
  MUX2_X1 M1_4_20 ( .A(\ML_int[4][20] ), .B(\ML_int[4][4] ), .S(n139), .Z(
        B[20]) );
  MUX2_X1 M1_4_19 ( .A(\ML_int[4][19] ), .B(\ML_int[4][3] ), .S(n139), .Z(
        B[19]) );
  MUX2_X1 M1_4_18 ( .A(\ML_int[4][18] ), .B(\ML_int[4][2] ), .S(n139), .Z(
        B[18]) );
  MUX2_X1 M1_4_17 ( .A(\ML_int[4][17] ), .B(\ML_int[4][1] ), .S(n139), .Z(
        B[17]) );
  MUX2_X1 M1_4_16 ( .A(\ML_int[4][16] ), .B(\ML_int[4][0] ), .S(n139), .Z(
        B[16]) );
  MUX2_X1 M0_4_15 ( .A(\ML_int[4][15] ), .B(\ML_int[4][31] ), .S(n139), .Z(
        B[15]) );
  MUX2_X1 M0_4_14 ( .A(\ML_int[4][14] ), .B(\ML_int[4][30] ), .S(n139), .Z(
        B[14]) );
  MUX2_X1 M0_4_13 ( .A(\ML_int[4][13] ), .B(\ML_int[4][29] ), .S(n138), .Z(
        B[13]) );
  MUX2_X1 M0_4_12 ( .A(\ML_int[4][12] ), .B(\ML_int[4][28] ), .S(n137), .Z(
        B[12]) );
  MUX2_X1 M0_4_11 ( .A(\ML_int[4][11] ), .B(\ML_int[4][27] ), .S(n137), .Z(
        B[11]) );
  MUX2_X1 M0_4_10 ( .A(\ML_int[4][10] ), .B(\ML_int[4][26] ), .S(n137), .Z(
        B[10]) );
  MUX2_X1 M0_4_9 ( .A(\ML_int[4][9] ), .B(\ML_int[4][25] ), .S(n137), .Z(B[9])
         );
  MUX2_X1 M0_4_8 ( .A(\ML_int[4][8] ), .B(\ML_int[4][24] ), .S(n137), .Z(B[8])
         );
  MUX2_X1 M0_4_7 ( .A(\ML_int[4][7] ), .B(\ML_int[4][23] ), .S(n137), .Z(B[7])
         );
  MUX2_X1 M0_4_6 ( .A(\ML_int[4][6] ), .B(\ML_int[4][22] ), .S(n137), .Z(B[6])
         );
  MUX2_X1 M0_4_5 ( .A(\ML_int[4][5] ), .B(\ML_int[4][21] ), .S(n137), .Z(B[5])
         );
  MUX2_X1 M0_4_4 ( .A(\ML_int[4][4] ), .B(\ML_int[4][20] ), .S(n137), .Z(B[4])
         );
  MUX2_X1 M0_4_3 ( .A(\ML_int[4][3] ), .B(\ML_int[4][19] ), .S(n137), .Z(B[3])
         );
  MUX2_X1 M0_4_2 ( .A(\ML_int[4][2] ), .B(\ML_int[4][18] ), .S(n137), .Z(B[2])
         );
  MUX2_X1 M0_4_1 ( .A(\ML_int[4][1] ), .B(\ML_int[4][17] ), .S(n137), .Z(B[1])
         );
  MUX2_X1 M0_4_0 ( .A(\ML_int[4][0] ), .B(\ML_int[4][16] ), .S(n139), .Z(B[0])
         );
  MUX2_X1 M1_3_31 ( .A(\ML_int[3][31] ), .B(\ML_int[3][23] ), .S(n135), .Z(
        \ML_int[4][31] ) );
  MUX2_X1 M1_3_30 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S(n135), .Z(
        \ML_int[4][30] ) );
  MUX2_X1 M1_3_29 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S(n135), .Z(
        \ML_int[4][29] ) );
  MUX2_X1 M1_3_28 ( .A(\ML_int[3][28] ), .B(\ML_int[3][20] ), .S(n135), .Z(
        \ML_int[4][28] ) );
  MUX2_X1 M1_3_27 ( .A(\ML_int[3][27] ), .B(\ML_int[3][19] ), .S(n135), .Z(
        \ML_int[4][27] ) );
  MUX2_X1 M1_3_26 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S(n135), .Z(
        \ML_int[4][26] ) );
  MUX2_X1 M1_3_25 ( .A(\ML_int[3][25] ), .B(\ML_int[3][17] ), .S(n135), .Z(
        \ML_int[4][25] ) );
  MUX2_X1 M1_3_24 ( .A(\ML_int[3][24] ), .B(\ML_int[3][16] ), .S(n134), .Z(
        \ML_int[4][24] ) );
  MUX2_X1 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S(n134), .Z(
        \ML_int[4][23] ) );
  MUX2_X1 M1_3_22 ( .A(\ML_int[3][22] ), .B(\ML_int[3][14] ), .S(n134), .Z(
        \ML_int[4][22] ) );
  MUX2_X1 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S(n134), .Z(
        \ML_int[4][21] ) );
  MUX2_X1 M1_3_20 ( .A(\ML_int[3][20] ), .B(\ML_int[3][12] ), .S(n136), .Z(
        \ML_int[4][20] ) );
  MUX2_X1 M1_3_19 ( .A(\ML_int[3][19] ), .B(\ML_int[3][11] ), .S(n134), .Z(
        \ML_int[4][19] ) );
  MUX2_X1 M1_3_18 ( .A(\ML_int[3][18] ), .B(\ML_int[3][10] ), .S(n135), .Z(
        \ML_int[4][18] ) );
  MUX2_X1 M1_3_17 ( .A(\ML_int[3][17] ), .B(\ML_int[3][9] ), .S(n136), .Z(
        \ML_int[4][17] ) );
  MUX2_X1 M1_3_16 ( .A(\ML_int[3][16] ), .B(\ML_int[3][8] ), .S(n136), .Z(
        \ML_int[4][16] ) );
  MUX2_X1 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S(n136), .Z(
        \ML_int[4][15] ) );
  MUX2_X1 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S(n136), .Z(
        \ML_int[4][14] ) );
  MUX2_X1 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S(n136), .Z(
        \ML_int[4][13] ) );
  MUX2_X1 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S(n136), .Z(
        \ML_int[4][12] ) );
  MUX2_X1 M1_3_11 ( .A(\ML_int[3][11] ), .B(\ML_int[3][3] ), .S(n136), .Z(
        \ML_int[4][11] ) );
  MUX2_X1 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S(n135), .Z(
        \ML_int[4][10] ) );
  MUX2_X1 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(n135), .Z(
        \ML_int[4][9] ) );
  MUX2_X1 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S(n135), .Z(
        \ML_int[4][8] ) );
  MUX2_X1 M0_3_7 ( .A(\ML_int[3][7] ), .B(\ML_int[3][31] ), .S(n135), .Z(
        \ML_int[4][7] ) );
  MUX2_X1 M0_3_6 ( .A(\ML_int[3][6] ), .B(\ML_int[3][30] ), .S(n134), .Z(
        \ML_int[4][6] ) );
  MUX2_X1 M0_3_5 ( .A(\ML_int[3][5] ), .B(\ML_int[3][29] ), .S(n134), .Z(
        \ML_int[4][5] ) );
  MUX2_X1 M0_3_4 ( .A(\ML_int[3][4] ), .B(\ML_int[3][28] ), .S(n134), .Z(
        \ML_int[4][4] ) );
  MUX2_X1 M0_3_3 ( .A(\ML_int[3][3] ), .B(\ML_int[3][27] ), .S(n134), .Z(
        \ML_int[4][3] ) );
  MUX2_X1 M0_3_2 ( .A(\ML_int[3][2] ), .B(\ML_int[3][26] ), .S(n134), .Z(
        \ML_int[4][2] ) );
  MUX2_X1 M0_3_1 ( .A(\ML_int[3][1] ), .B(\ML_int[3][25] ), .S(n134), .Z(
        \ML_int[4][1] ) );
  MUX2_X1 M0_3_0 ( .A(\ML_int[3][0] ), .B(\ML_int[3][24] ), .S(n134), .Z(
        \ML_int[4][0] ) );
  MUX2_X1 M1_2_31 ( .A(\ML_int[2][31] ), .B(\ML_int[2][27] ), .S(n133), .Z(
        \ML_int[3][31] ) );
  MUX2_X1 M1_2_30 ( .A(\ML_int[2][30] ), .B(\ML_int[2][26] ), .S(n132), .Z(
        \ML_int[3][30] ) );
  MUX2_X1 M1_2_29 ( .A(\ML_int[2][29] ), .B(\ML_int[2][25] ), .S(n132), .Z(
        \ML_int[3][29] ) );
  MUX2_X1 M1_2_28 ( .A(\ML_int[2][28] ), .B(\ML_int[2][24] ), .S(n132), .Z(
        \ML_int[3][28] ) );
  MUX2_X1 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(n132), .Z(
        \ML_int[3][27] ) );
  MUX2_X1 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(n132), .Z(
        \ML_int[3][26] ) );
  MUX2_X1 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(n132), .Z(
        \ML_int[3][25] ) );
  MUX2_X1 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(n132), .Z(
        \ML_int[3][24] ) );
  MUX2_X1 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(n132), .Z(
        \ML_int[3][23] ) );
  MUX2_X1 M1_2_22 ( .A(\ML_int[2][22] ), .B(\ML_int[2][18] ), .S(n132), .Z(
        \ML_int[3][22] ) );
  MUX2_X1 M1_2_21 ( .A(\ML_int[2][21] ), .B(\ML_int[2][17] ), .S(n132), .Z(
        \ML_int[3][21] ) );
  MUX2_X1 M1_2_20 ( .A(\ML_int[2][20] ), .B(\ML_int[2][16] ), .S(n132), .Z(
        \ML_int[3][20] ) );
  MUX2_X1 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S(n132), .Z(
        \ML_int[3][19] ) );
  MUX2_X1 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(n131), .Z(
        \ML_int[3][18] ) );
  MUX2_X1 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(n133), .Z(
        \ML_int[3][17] ) );
  MUX2_X1 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S(n133), .Z(
        \ML_int[3][16] ) );
  MUX2_X1 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S(n133), .Z(
        \ML_int[3][15] ) );
  MUX2_X1 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S(n133), .Z(
        \ML_int[3][14] ) );
  MUX2_X1 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S(n133), .Z(
        \ML_int[3][13] ) );
  MUX2_X1 M1_2_12 ( .A(\ML_int[2][12] ), .B(\ML_int[2][8] ), .S(n133), .Z(
        \ML_int[3][12] ) );
  MUX2_X1 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(n133), .Z(
        \ML_int[3][11] ) );
  MUX2_X1 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(n131), .Z(
        \ML_int[3][10] ) );
  MUX2_X1 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(n131), .Z(
        \ML_int[3][9] ) );
  MUX2_X1 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(n131), .Z(
        \ML_int[3][8] ) );
  MUX2_X1 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(n131), .Z(
        \ML_int[3][7] ) );
  MUX2_X1 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(n131), .Z(
        \ML_int[3][6] ) );
  MUX2_X1 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S(n131), .Z(
        \ML_int[3][5] ) );
  MUX2_X1 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(n131), .Z(
        \ML_int[3][4] ) );
  MUX2_X1 M0_2_3 ( .A(\ML_int[2][3] ), .B(\ML_int[2][31] ), .S(n131), .Z(
        \ML_int[3][3] ) );
  MUX2_X1 M0_2_2 ( .A(\ML_int[2][2] ), .B(\ML_int[2][30] ), .S(n131), .Z(
        \ML_int[3][2] ) );
  MUX2_X1 M0_2_1 ( .A(\ML_int[2][1] ), .B(\ML_int[2][29] ), .S(n131), .Z(
        \ML_int[3][1] ) );
  MUX2_X1 M0_2_0 ( .A(\ML_int[2][0] ), .B(\ML_int[2][28] ), .S(n131), .Z(
        \ML_int[3][0] ) );
  MUX2_X1 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(n129), .Z(
        \ML_int[2][31] ) );
  MUX2_X1 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S(n129), .Z(
        \ML_int[2][30] ) );
  MUX2_X1 M1_1_29 ( .A(\ML_int[1][29] ), .B(\ML_int[1][27] ), .S(n129), .Z(
        \ML_int[2][29] ) );
  MUX2_X1 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S(n129), .Z(
        \ML_int[2][28] ) );
  MUX2_X1 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S(n129), .Z(
        \ML_int[2][27] ) );
  MUX2_X1 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S(n129), .Z(
        \ML_int[2][26] ) );
  MUX2_X1 M1_1_25 ( .A(\ML_int[1][25] ), .B(\ML_int[1][23] ), .S(n129), .Z(
        \ML_int[2][25] ) );
  MUX2_X1 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(n128), .Z(
        \ML_int[2][24] ) );
  MUX2_X1 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S(n128), .Z(
        \ML_int[2][23] ) );
  MUX2_X1 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(n128), .Z(
        \ML_int[2][22] ) );
  MUX2_X1 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(n128), .Z(
        \ML_int[2][21] ) );
  MUX2_X1 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S(n128), .Z(
        \ML_int[2][20] ) );
  MUX2_X1 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(n128), .Z(
        \ML_int[2][19] ) );
  MUX2_X1 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S(n128), .Z(
        \ML_int[2][18] ) );
  MUX2_X1 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S(n130), .Z(
        \ML_int[2][17] ) );
  MUX2_X1 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(n130), .Z(
        \ML_int[2][16] ) );
  MUX2_X1 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(n130), .Z(
        \ML_int[2][15] ) );
  MUX2_X1 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S(n130), .Z(
        \ML_int[2][14] ) );
  MUX2_X1 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(n130), .Z(
        \ML_int[2][13] ) );
  MUX2_X1 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S(n130), .Z(
        \ML_int[2][12] ) );
  MUX2_X1 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(n130), .Z(
        \ML_int[2][11] ) );
  MUX2_X1 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(n129), .Z(
        \ML_int[2][10] ) );
  MUX2_X1 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(n128), .Z(
        \ML_int[2][9] ) );
  MUX2_X1 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(n129), .Z(
        \ML_int[2][8] ) );
  MUX2_X1 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(n128), .Z(
        \ML_int[2][7] ) );
  MUX2_X1 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(n128), .Z(
        \ML_int[2][6] ) );
  MUX2_X1 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(n128), .Z(
        \ML_int[2][5] ) );
  MUX2_X1 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(n129), .Z(
        \ML_int[2][4] ) );
  MUX2_X1 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(n130), .Z(
        \ML_int[2][3] ) );
  MUX2_X1 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(n129), .Z(
        \ML_int[2][2] ) );
  MUX2_X1 M0_1_1 ( .A(\ML_int[1][1] ), .B(\ML_int[1][31] ), .S(n129), .Z(
        \ML_int[2][1] ) );
  MUX2_X1 M0_1_0 ( .A(\ML_int[1][0] ), .B(\ML_int[1][30] ), .S(n128), .Z(
        \ML_int[2][0] ) );
  MUX2_X1 M1_0_31 ( .A(A[31]), .B(A[30]), .S(n126), .Z(\ML_int[1][31] ) );
  MUX2_X1 M1_0_30 ( .A(A[30]), .B(A[29]), .S(n126), .Z(\ML_int[1][30] ) );
  MUX2_X1 M1_0_29 ( .A(A[29]), .B(A[28]), .S(n126), .Z(\ML_int[1][29] ) );
  MUX2_X1 M1_0_28 ( .A(A[28]), .B(A[27]), .S(n126), .Z(\ML_int[1][28] ) );
  MUX2_X1 M1_0_27 ( .A(A[27]), .B(A[26]), .S(n126), .Z(\ML_int[1][27] ) );
  MUX2_X1 M1_0_26 ( .A(A[26]), .B(A[25]), .S(n126), .Z(\ML_int[1][26] ) );
  MUX2_X1 M1_0_25 ( .A(A[25]), .B(A[24]), .S(n126), .Z(\ML_int[1][25] ) );
  MUX2_X1 M1_0_24 ( .A(A[24]), .B(A[23]), .S(n126), .Z(\ML_int[1][24] ) );
  MUX2_X1 M1_0_23 ( .A(A[23]), .B(A[22]), .S(n126), .Z(\ML_int[1][23] ) );
  MUX2_X1 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n125), .Z(\ML_int[1][22] ) );
  MUX2_X1 M1_0_21 ( .A(A[21]), .B(A[20]), .S(n125), .Z(\ML_int[1][21] ) );
  MUX2_X1 M1_0_20 ( .A(A[20]), .B(A[19]), .S(n126), .Z(\ML_int[1][20] ) );
  MUX2_X1 M1_0_19 ( .A(A[19]), .B(A[18]), .S(n126), .Z(\ML_int[1][19] ) );
  MUX2_X1 M1_0_18 ( .A(A[18]), .B(A[17]), .S(n125), .Z(\ML_int[1][18] ) );
  MUX2_X1 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n125), .Z(\ML_int[1][17] ) );
  MUX2_X1 M1_0_16 ( .A(A[16]), .B(A[15]), .S(n125), .Z(\ML_int[1][16] ) );
  MUX2_X1 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n125), .Z(\ML_int[1][15] ) );
  MUX2_X1 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n125), .Z(\ML_int[1][14] ) );
  MUX2_X1 M1_0_13 ( .A(A[13]), .B(A[12]), .S(n125), .Z(\ML_int[1][13] ) );
  MUX2_X1 M1_0_12 ( .A(A[12]), .B(A[11]), .S(n125), .Z(\ML_int[1][12] ) );
  MUX2_X1 M1_0_11 ( .A(A[11]), .B(A[10]), .S(n125), .Z(\ML_int[1][11] ) );
  MUX2_X1 M1_0_10 ( .A(A[10]), .B(A[9]), .S(n127), .Z(\ML_int[1][10] ) );
  MUX2_X1 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n127), .Z(\ML_int[1][9] ) );
  MUX2_X1 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n127), .Z(\ML_int[1][8] ) );
  MUX2_X1 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n127), .Z(\ML_int[1][7] ) );
  MUX2_X1 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n127), .Z(\ML_int[1][6] ) );
  MUX2_X1 M1_0_5 ( .A(A[5]), .B(A[4]), .S(n126), .Z(\ML_int[1][5] ) );
  MUX2_X1 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n125), .Z(\ML_int[1][4] ) );
  MUX2_X1 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n127), .Z(\ML_int[1][3] ) );
  MUX2_X1 M1_0_2 ( .A(A[2]), .B(A[1]), .S(n127), .Z(\ML_int[1][2] ) );
  MUX2_X1 M1_0_1 ( .A(A[1]), .B(A[0]), .S(n127), .Z(\ML_int[1][1] ) );
  MUX2_X1 M0_0_0 ( .A(A[0]), .B(A[31]), .S(n125), .Z(\ML_int[1][0] ) );
  BUF_X1 U2 ( .A(SH[1]), .Z(n128) );
  BUF_X1 U3 ( .A(SH[1]), .Z(n129) );
  BUF_X1 U4 ( .A(SH[3]), .Z(n134) );
  BUF_X1 U5 ( .A(SH[3]), .Z(n135) );
  BUF_X1 U6 ( .A(SH[4]), .Z(n137) );
  BUF_X1 U7 ( .A(SH[4]), .Z(n138) );
  BUF_X1 U8 ( .A(SH[1]), .Z(n130) );
  BUF_X1 U9 ( .A(SH[3]), .Z(n136) );
  BUF_X1 U10 ( .A(SH[4]), .Z(n139) );
  BUF_X1 U11 ( .A(SH[0]), .Z(n125) );
  BUF_X1 U12 ( .A(SH[0]), .Z(n126) );
  BUF_X1 U13 ( .A(SH[2]), .Z(n131) );
  BUF_X1 U14 ( .A(SH[2]), .Z(n132) );
  BUF_X1 U15 ( .A(SH[0]), .Z(n127) );
  BUF_X1 U16 ( .A(SH[2]), .Z(n133) );
endmodule


module SHIFTER_GENERIC_N32_DW_sra_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \A[31] , n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355;
  assign B[31] = \A[31] ;
  assign \A[31]  = A[31];

  NOR2_X2 U2 ( .A1(SH[2]), .A2(SH[3]), .ZN(n104) );
  MUX2_X1 U174 ( .A(\A[31] ), .B(A[30]), .S(n86), .Z(n115) );
  NAND2_X1 U3 ( .A1(n342), .A2(\A[31] ), .ZN(n91) );
  INV_X1 U4 ( .A(n75), .ZN(n43) );
  INV_X1 U5 ( .A(n342), .ZN(n338) );
  INV_X1 U6 ( .A(n88), .ZN(n83) );
  INV_X1 U7 ( .A(n85), .ZN(n80) );
  OAI221_X1 U8 ( .B1(n63), .B2(n40), .C1(n64), .C2(n338), .A(n65), .ZN(B[6])
         );
  OAI221_X1 U9 ( .B1(n50), .B2(n40), .C1(n51), .C2(n338), .A(n52), .ZN(B[8])
         );
  OAI221_X1 U10 ( .B1(n39), .B2(n40), .C1(n41), .C2(n338), .A(n42), .ZN(B[9])
         );
  OAI221_X1 U11 ( .B1(n150), .B2(n40), .C1(n98), .C2(n338), .A(n151), .ZN(
        B[12]) );
  OAI221_X1 U12 ( .B1(n143), .B2(n40), .C1(n97), .C2(n338), .A(n144), .ZN(
        B[13]) );
  NAND2_X1 U13 ( .A1(n102), .A2(n338), .ZN(n75) );
  INV_X1 U14 ( .A(n40), .ZN(n78) );
  BUF_X1 U15 ( .A(n336), .Z(n339) );
  BUF_X1 U16 ( .A(n336), .Z(n340) );
  BUF_X1 U17 ( .A(n337), .Z(n341) );
  BUF_X1 U18 ( .A(n337), .Z(n342) );
  NOR2_X1 U19 ( .A1(n335), .A2(SH[3]), .ZN(n102) );
  INV_X1 U20 ( .A(n89), .ZN(n84) );
  NOR2_X1 U21 ( .A1(n334), .A2(SH[1]), .ZN(n85) );
  INV_X1 U22 ( .A(n86), .ZN(n81) );
  NAND2_X1 U23 ( .A1(n104), .A2(n338), .ZN(n40) );
  AOI221_X1 U24 ( .B1(n85), .B2(A[7]), .C1(n86), .C2(A[6]), .A(n96), .ZN(n63)
         );
  OAI22_X1 U25 ( .A1(n349), .A2(n88), .B1(n350), .B2(n89), .ZN(n96) );
  AOI221_X1 U26 ( .B1(n108), .B2(n102), .C1(n109), .C2(n104), .A(n105), .ZN(
        n58) );
  AOI221_X1 U27 ( .B1(n106), .B2(n102), .C1(n107), .C2(n104), .A(n105), .ZN(
        n51) );
  AOI221_X1 U28 ( .B1(n101), .B2(n102), .C1(n103), .C2(n104), .A(n105), .ZN(
        n41) );
  AOI221_X1 U29 ( .B1(n115), .B2(n102), .C1(n110), .C2(n104), .A(n105), .ZN(
        n100) );
  AOI221_X1 U30 ( .B1(n55), .B2(n102), .C1(n54), .C2(n104), .A(n173), .ZN(n135) );
  INV_X1 U31 ( .A(n174), .ZN(n173) );
  AOI22_X1 U32 ( .A1(n132), .A2(n106), .B1(n114), .B2(n107), .ZN(n174) );
  AOI221_X1 U33 ( .B1(n48), .B2(n102), .C1(n46), .C2(n104), .A(n133), .ZN(n121) );
  INV_X1 U34 ( .A(n134), .ZN(n133) );
  AOI22_X1 U35 ( .A1(n132), .A2(n101), .B1(n114), .B2(n103), .ZN(n134) );
  AOI221_X1 U36 ( .B1(n111), .B2(n102), .C1(n68), .C2(n104), .A(n130), .ZN(n92) );
  INV_X1 U37 ( .A(n131), .ZN(n130) );
  AOI22_X1 U38 ( .A1(n132), .A2(n115), .B1(n114), .B2(n110), .ZN(n131) );
  AOI221_X1 U39 ( .B1(n109), .B2(n102), .C1(n62), .C2(n104), .A(n127), .ZN(n76) );
  INV_X1 U40 ( .A(n128), .ZN(n127) );
  AOI21_X1 U41 ( .B1(n114), .B2(n108), .A(n116), .ZN(n128) );
  AOI221_X1 U42 ( .B1(n107), .B2(n102), .C1(n55), .C2(n104), .A(n119), .ZN(n73) );
  INV_X1 U43 ( .A(n120), .ZN(n119) );
  AOI21_X1 U44 ( .B1(n114), .B2(n106), .A(n116), .ZN(n120) );
  AOI221_X1 U45 ( .B1(n103), .B2(n102), .C1(n48), .C2(n104), .A(n117), .ZN(n70) );
  INV_X1 U46 ( .A(n118), .ZN(n117) );
  AOI21_X1 U47 ( .B1(n114), .B2(n101), .A(n116), .ZN(n118) );
  AOI221_X1 U48 ( .B1(n110), .B2(n102), .C1(n111), .C2(n104), .A(n112), .ZN(
        n64) );
  INV_X1 U49 ( .A(n113), .ZN(n112) );
  AOI21_X1 U50 ( .B1(n114), .B2(n115), .A(n116), .ZN(n113) );
  AOI222_X1 U51 ( .A1(n43), .A2(n61), .B1(n45), .B2(n62), .C1(n47), .C2(n109), 
        .ZN(n153) );
  AOI222_X1 U52 ( .A1(n43), .A2(n67), .B1(n45), .B2(n68), .C1(n47), .C2(n111), 
        .ZN(n160) );
  AOI222_X1 U53 ( .A1(n43), .A2(n54), .B1(n45), .B2(n55), .C1(n47), .C2(n107), 
        .ZN(n151) );
  AOI222_X1 U54 ( .A1(n43), .A2(n66), .B1(n45), .B2(n67), .C1(n47), .C2(n68), 
        .ZN(n65) );
  AOI222_X1 U55 ( .A1(n43), .A2(n60), .B1(n45), .B2(n61), .C1(n47), .C2(n62), 
        .ZN(n59) );
  AOI222_X1 U56 ( .A1(n43), .A2(n53), .B1(n45), .B2(n54), .C1(n47), .C2(n55), 
        .ZN(n52) );
  AOI222_X1 U57 ( .A1(n43), .A2(n56), .B1(n45), .B2(n53), .C1(n47), .C2(n54), 
        .ZN(n74) );
  AOI222_X1 U58 ( .A1(n43), .A2(n49), .B1(n45), .B2(n44), .C1(n47), .C2(n46), 
        .ZN(n71) );
  AOI222_X1 U59 ( .A1(n43), .A2(n44), .B1(n45), .B2(n46), .C1(n47), .C2(n48), 
        .ZN(n42) );
  AOI222_X1 U60 ( .A1(n43), .A2(n46), .B1(n45), .B2(n48), .C1(n47), .C2(n103), 
        .ZN(n144) );
  AOI222_X1 U61 ( .A1(n43), .A2(n68), .B1(n45), .B2(n111), .C1(n47), .C2(n110), 
        .ZN(n141) );
  OAI221_X1 U62 ( .B1(n57), .B2(n75), .C1(n76), .C2(n338), .A(n77), .ZN(B[3])
         );
  OAI221_X1 U63 ( .B1(n72), .B2(n40), .C1(n73), .C2(n338), .A(n74), .ZN(B[4])
         );
  OAI221_X1 U64 ( .B1(n69), .B2(n40), .C1(n70), .C2(n338), .A(n71), .ZN(B[5])
         );
  OAI221_X1 U65 ( .B1(n57), .B2(n40), .C1(n58), .C2(n338), .A(n59), .ZN(B[7])
         );
  OAI221_X1 U66 ( .B1(n72), .B2(n75), .C1(n135), .C2(n338), .A(n167), .ZN(B[0]) );
  OAI221_X1 U67 ( .B1(n69), .B2(n75), .C1(n121), .C2(n338), .A(n122), .ZN(B[1]) );
  OAI221_X1 U68 ( .B1(n63), .B2(n75), .C1(n92), .C2(n338), .A(n93), .ZN(B[2])
         );
  OAI221_X1 U69 ( .B1(n159), .B2(n40), .C1(n100), .C2(n338), .A(n160), .ZN(
        B[10]) );
  OAI221_X1 U70 ( .B1(n152), .B2(n40), .C1(n99), .C2(n338), .A(n153), .ZN(
        B[11]) );
  OAI221_X1 U71 ( .B1(n140), .B2(n40), .C1(n90), .C2(n338), .A(n141), .ZN(
        B[14]) );
  OAI221_X1 U72 ( .B1(n136), .B2(n75), .C1(n137), .C2(n40), .A(n138), .ZN(
        B[15]) );
  OAI21_X1 U73 ( .B1(n339), .B2(n135), .A(n91), .ZN(B[16]) );
  OAI21_X1 U74 ( .B1(n339), .B2(n121), .A(n91), .ZN(B[17]) );
  OAI21_X1 U75 ( .B1(n339), .B2(n92), .A(n91), .ZN(B[18]) );
  OAI21_X1 U76 ( .B1(n339), .B2(n76), .A(n91), .ZN(B[19]) );
  OAI21_X1 U77 ( .B1(n340), .B2(n73), .A(n91), .ZN(B[20]) );
  OAI21_X1 U78 ( .B1(n340), .B2(n70), .A(n91), .ZN(B[21]) );
  OAI21_X1 U79 ( .B1(n340), .B2(n64), .A(n91), .ZN(B[22]) );
  OAI21_X1 U80 ( .B1(n340), .B2(n58), .A(n91), .ZN(B[23]) );
  OAI21_X1 U81 ( .B1(n339), .B2(n51), .A(n91), .ZN(B[24]) );
  OAI21_X1 U82 ( .B1(n340), .B2(n41), .A(n91), .ZN(B[25]) );
  OAI21_X1 U83 ( .B1(n341), .B2(n100), .A(n91), .ZN(B[26]) );
  OAI21_X1 U84 ( .B1(n341), .B2(n99), .A(n91), .ZN(B[27]) );
  OAI21_X1 U85 ( .B1(n341), .B2(n98), .A(n91), .ZN(B[28]) );
  OAI21_X1 U86 ( .B1(n341), .B2(n97), .A(n91), .ZN(B[29]) );
  OAI21_X1 U87 ( .B1(n341), .B2(n90), .A(n91), .ZN(B[30]) );
  AOI221_X1 U88 ( .B1(n47), .B2(n108), .C1(n45), .C2(n109), .A(n139), .ZN(n138) );
  INV_X1 U89 ( .A(n91), .ZN(n139) );
  NAND2_X1 U90 ( .A1(SH[1]), .A2(n334), .ZN(n88) );
  NOR2_X1 U91 ( .A1(n129), .A2(n335), .ZN(n116) );
  AND2_X1 U92 ( .A1(n170), .A2(n335), .ZN(n45) );
  AND2_X1 U93 ( .A1(SH[3]), .A2(n335), .ZN(n114) );
  AOI21_X1 U94 ( .B1(n108), .B2(n104), .A(n142), .ZN(n99) );
  AOI21_X1 U95 ( .B1(n106), .B2(n104), .A(n142), .ZN(n98) );
  AOI21_X1 U96 ( .B1(n101), .B2(n104), .A(n142), .ZN(n97) );
  AOI21_X1 U97 ( .B1(n115), .B2(n104), .A(n142), .ZN(n90) );
  INV_X1 U98 ( .A(n129), .ZN(n105) );
  INV_X1 U99 ( .A(n140), .ZN(n67) );
  INV_X1 U100 ( .A(n137), .ZN(n61) );
  INV_X1 U101 ( .A(n62), .ZN(n136) );
  INV_X1 U102 ( .A(n53), .ZN(n150) );
  INV_X1 U103 ( .A(n44), .ZN(n143) );
  AND2_X1 U104 ( .A1(SH[3]), .A2(n338), .ZN(n170) );
  INV_X1 U105 ( .A(n56), .ZN(n50) );
  INV_X1 U106 ( .A(n49), .ZN(n39) );
  INV_X1 U107 ( .A(n66), .ZN(n159) );
  INV_X1 U108 ( .A(n60), .ZN(n152) );
  BUF_X1 U109 ( .A(SH[4]), .Z(n337) );
  BUF_X1 U110 ( .A(SH[4]), .Z(n336) );
  NOR2_X1 U111 ( .A1(SH[0]), .A2(SH[1]), .ZN(n86) );
  OAI221_X1 U112 ( .B1(n80), .B2(n37), .C1(n81), .C2(n36), .A(n176), .ZN(n106)
         );
  INV_X1 U113 ( .A(A[29]), .ZN(n37) );
  AOI22_X1 U114 ( .A1(A[30]), .A2(n83), .B1(\A[31] ), .B2(n84), .ZN(n176) );
  OAI221_X1 U115 ( .B1(n80), .B2(n32), .C1(n81), .C2(n31), .A(n154), .ZN(n109)
         );
  AOI22_X1 U116 ( .A1(A[25]), .A2(n83), .B1(A[26]), .B2(n84), .ZN(n154) );
  OAI221_X1 U117 ( .B1(n80), .B2(n33), .C1(n81), .C2(n32), .A(n175), .ZN(n107)
         );
  AOI22_X1 U118 ( .A1(A[26]), .A2(n83), .B1(A[27]), .B2(n84), .ZN(n175) );
  OAI221_X1 U119 ( .B1(n80), .B2(n34), .C1(n81), .C2(n33), .A(n145), .ZN(n103)
         );
  AOI22_X1 U120 ( .A1(A[27]), .A2(n83), .B1(A[28]), .B2(n84), .ZN(n145) );
  OAI221_X1 U121 ( .B1(n80), .B2(n35), .C1(n81), .C2(n34), .A(n165), .ZN(n110)
         );
  AOI22_X1 U122 ( .A1(A[28]), .A2(n83), .B1(A[29]), .B2(n84), .ZN(n165) );
  OAI221_X1 U123 ( .B1(n80), .B2(n29), .C1(n28), .C2(n81), .A(n178), .ZN(n55)
         );
  AOI22_X1 U124 ( .A1(A[22]), .A2(n83), .B1(A[23]), .B2(n84), .ZN(n178) );
  OAI221_X1 U125 ( .B1(n80), .B2(n30), .C1(n81), .C2(n29), .A(n146), .ZN(n48)
         );
  AOI22_X1 U126 ( .A1(A[23]), .A2(n83), .B1(A[24]), .B2(n84), .ZN(n146) );
  OAI221_X1 U127 ( .B1(n80), .B2(n31), .C1(n81), .C2(n30), .A(n161), .ZN(n111)
         );
  AOI22_X1 U128 ( .A1(A[24]), .A2(n83), .B1(A[25]), .B2(n84), .ZN(n161) );
  OAI221_X1 U129 ( .B1(n80), .B2(n354), .C1(n81), .C2(n353), .A(n172), .ZN(n53) );
  AOI22_X1 U130 ( .A1(A[14]), .A2(n83), .B1(A[15]), .B2(n84), .ZN(n172) );
  OAI221_X1 U131 ( .B1(n80), .B2(n355), .C1(n81), .C2(n354), .A(n149), .ZN(n44) );
  AOI22_X1 U132 ( .A1(A[15]), .A2(n83), .B1(A[16]), .B2(n84), .ZN(n149) );
  OAI221_X1 U133 ( .B1(n80), .B2(n26), .C1(n81), .C2(n25), .A(n147), .ZN(n46)
         );
  AOI22_X1 U134 ( .A1(A[19]), .A2(n83), .B1(A[20]), .B2(n84), .ZN(n147) );
  OAI221_X1 U135 ( .B1(n80), .B2(n36), .C1(n81), .C2(n35), .A(n157), .ZN(n108)
         );
  AOI22_X1 U136 ( .A1(A[29]), .A2(n83), .B1(A[30]), .B2(n84), .ZN(n157) );
  OAI221_X1 U137 ( .B1(n28), .B2(n80), .C1(n27), .C2(n81), .A(n155), .ZN(n62)
         );
  AOI22_X1 U138 ( .A1(A[21]), .A2(n83), .B1(A[22]), .B2(n84), .ZN(n155) );
  OAI221_X1 U139 ( .B1(n27), .B2(n80), .C1(n26), .C2(n81), .A(n162), .ZN(n68)
         );
  AOI22_X1 U140 ( .A1(A[20]), .A2(n83), .B1(A[21]), .B2(n84), .ZN(n162) );
  OAI221_X1 U141 ( .B1(n88), .B2(n26), .C1(n27), .C2(n89), .A(n177), .ZN(n54)
         );
  AOI22_X1 U142 ( .A1(A[17]), .A2(n85), .B1(A[16]), .B2(n86), .ZN(n177) );
  AOI221_X1 U143 ( .B1(n85), .B2(A[5]), .C1(n86), .C2(A[4]), .A(n179), .ZN(n72) );
  OAI22_X1 U144 ( .A1(n347), .A2(n88), .B1(n348), .B2(n89), .ZN(n179) );
  AOI221_X1 U145 ( .B1(n85), .B2(A[8]), .C1(n86), .C2(A[7]), .A(n87), .ZN(n57)
         );
  OAI22_X1 U146 ( .A1(n350), .A2(n88), .B1(n351), .B2(n89), .ZN(n87) );
  AOI221_X1 U147 ( .B1(n85), .B2(A[6]), .C1(n86), .C2(A[5]), .A(n126), .ZN(n69) );
  OAI22_X1 U148 ( .A1(n348), .A2(n88), .B1(n349), .B2(n89), .ZN(n126) );
  AOI221_X1 U149 ( .B1(n85), .B2(A[15]), .C1(n86), .C2(A[14]), .A(n163), .ZN(
        n140) );
  INV_X1 U150 ( .A(n164), .ZN(n163) );
  AOI22_X1 U151 ( .A1(A[16]), .A2(n83), .B1(A[17]), .B2(n84), .ZN(n164) );
  OAI221_X1 U152 ( .B1(n80), .B2(n350), .C1(n81), .C2(n349), .A(n169), .ZN(n56) );
  AOI22_X1 U153 ( .A1(A[10]), .A2(n83), .B1(A[11]), .B2(n84), .ZN(n169) );
  OAI221_X1 U154 ( .B1(n80), .B2(n351), .C1(n81), .C2(n350), .A(n124), .ZN(n49) );
  AOI22_X1 U155 ( .A1(A[11]), .A2(n83), .B1(A[12]), .B2(n84), .ZN(n124) );
  OAI221_X1 U156 ( .B1(n80), .B2(n352), .C1(n81), .C2(n351), .A(n166), .ZN(n66) );
  AOI22_X1 U157 ( .A1(A[12]), .A2(n83), .B1(A[13]), .B2(n84), .ZN(n166) );
  OAI221_X1 U158 ( .B1(n80), .B2(n353), .C1(n81), .C2(n352), .A(n158), .ZN(n60) );
  AOI22_X1 U159 ( .A1(A[13]), .A2(n83), .B1(A[14]), .B2(n84), .ZN(n158) );
  AOI221_X1 U160 ( .B1(n85), .B2(A[16]), .C1(n86), .C2(A[15]), .A(n156), .ZN(
        n137) );
  OAI22_X1 U161 ( .A1(n25), .A2(n88), .B1(n26), .B2(n89), .ZN(n156) );
  AOI222_X1 U162 ( .A1(n47), .A2(n44), .B1(n78), .B2(n123), .C1(n45), .C2(n49), 
        .ZN(n122) );
  OAI221_X1 U163 ( .B1(n80), .B2(n344), .C1(n81), .C2(n343), .A(n125), .ZN(
        n123) );
  AOI22_X1 U164 ( .A1(A[3]), .A2(n83), .B1(A[4]), .B2(n84), .ZN(n125) );
  AOI222_X1 U165 ( .A1(n47), .A2(n67), .B1(n78), .B2(n94), .C1(n45), .C2(n66), 
        .ZN(n93) );
  OAI221_X1 U166 ( .B1(n80), .B2(n345), .C1(n81), .C2(n344), .A(n95), .ZN(n94)
         );
  AOI22_X1 U167 ( .A1(A[4]), .A2(n83), .B1(A[5]), .B2(n84), .ZN(n95) );
  AOI222_X1 U168 ( .A1(n47), .A2(n61), .B1(n78), .B2(n79), .C1(n45), .C2(n60), 
        .ZN(n77) );
  OAI221_X1 U169 ( .B1(n80), .B2(n346), .C1(n81), .C2(n345), .A(n82), .ZN(n79)
         );
  AOI22_X1 U170 ( .A1(A[5]), .A2(n83), .B1(A[6]), .B2(n84), .ZN(n82) );
  AOI222_X1 U171 ( .A1(n47), .A2(n53), .B1(n78), .B2(n168), .C1(n45), .C2(n56), 
        .ZN(n167) );
  OAI221_X1 U172 ( .B1(n88), .B2(n344), .C1(n89), .C2(n345), .A(n171), .ZN(
        n168) );
  AOI22_X1 U173 ( .A1(A[1]), .A2(n85), .B1(A[0]), .B2(n86), .ZN(n171) );
  OAI21_X1 U175 ( .B1(n335), .B2(n38), .A(n129), .ZN(n142) );
  INV_X1 U176 ( .A(\A[31] ), .ZN(n38) );
  NAND2_X1 U177 ( .A1(SH[0]), .A2(SH[1]), .ZN(n89) );
  AND2_X1 U178 ( .A1(SH[2]), .A2(n170), .ZN(n47) );
  NAND2_X1 U179 ( .A1(\A[31] ), .A2(SH[3]), .ZN(n129) );
  INV_X1 U180 ( .A(n148), .ZN(n101) );
  AOI222_X1 U181 ( .A1(n86), .A2(A[29]), .B1(n85), .B2(A[30]), .C1(SH[1]), 
        .C2(\A[31] ), .ZN(n148) );
  INV_X1 U182 ( .A(A[18]), .ZN(n26) );
  AND2_X1 U183 ( .A1(SH[2]), .A2(SH[3]), .ZN(n132) );
  INV_X1 U184 ( .A(A[19]), .ZN(n27) );
  INV_X1 U185 ( .A(A[7]), .ZN(n348) );
  INV_X1 U186 ( .A(A[20]), .ZN(n28) );
  INV_X1 U187 ( .A(A[17]), .ZN(n25) );
  INV_X1 U188 ( .A(A[25]), .ZN(n33) );
  INV_X1 U189 ( .A(A[21]), .ZN(n29) );
  INV_X1 U190 ( .A(A[26]), .ZN(n34) );
  INV_X1 U191 ( .A(A[22]), .ZN(n30) );
  INV_X1 U192 ( .A(A[23]), .ZN(n31) );
  INV_X1 U193 ( .A(A[24]), .ZN(n32) );
  INV_X1 U194 ( .A(A[27]), .ZN(n35) );
  INV_X1 U195 ( .A(A[28]), .ZN(n36) );
  INV_X1 U196 ( .A(SH[0]), .ZN(n334) );
  INV_X1 U197 ( .A(SH[2]), .ZN(n335) );
  INV_X1 U198 ( .A(A[1]), .ZN(n343) );
  INV_X1 U199 ( .A(A[2]), .ZN(n344) );
  INV_X1 U200 ( .A(A[3]), .ZN(n345) );
  INV_X1 U201 ( .A(A[4]), .ZN(n346) );
  INV_X1 U202 ( .A(A[6]), .ZN(n347) );
  INV_X1 U203 ( .A(A[8]), .ZN(n349) );
  INV_X1 U204 ( .A(A[9]), .ZN(n350) );
  INV_X1 U205 ( .A(A[10]), .ZN(n351) );
  INV_X1 U206 ( .A(A[11]), .ZN(n352) );
  INV_X1 U207 ( .A(A[12]), .ZN(n353) );
  INV_X1 U208 ( .A(A[13]), .ZN(n354) );
  INV_X1 U209 ( .A(A[14]), .ZN(n355) );
endmodule


module SHIFTER_GENERIC_N32_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362;

  NOR2_X2 U5 ( .A1(SH[0]), .A2(SH[1]), .ZN(n84) );
  NOR2_X2 U6 ( .A1(n339), .A2(SH[1]), .ZN(n83) );
  MUX2_X1 U137 ( .A(n106), .B(n90), .S(SH[2]), .Z(n117) );
  NOR2_X1 U3 ( .A1(n340), .A2(n341), .ZN(n104) );
  INV_X1 U4 ( .A(n39), .ZN(n77) );
  NAND2_X1 U7 ( .A1(n103), .A2(n349), .ZN(n39) );
  INV_X1 U8 ( .A(n346), .ZN(n349) );
  INV_X1 U9 ( .A(n169), .ZN(n86) );
  INV_X1 U10 ( .A(n74), .ZN(n42) );
  INV_X1 U11 ( .A(n83), .ZN(n88) );
  OAI221_X1 U12 ( .B1(n60), .B2(n39), .C1(n61), .C2(n349), .A(n62), .ZN(B[6])
         );
  OAI221_X1 U13 ( .B1(n48), .B2(n39), .C1(n49), .C2(n349), .A(n50), .ZN(B[8])
         );
  OAI221_X1 U14 ( .B1(n38), .B2(n39), .C1(n40), .C2(n349), .A(n41), .ZN(B[9])
         );
  INV_X1 U15 ( .A(n138), .ZN(B[12]) );
  OAI221_X1 U16 ( .B1(n131), .B2(n74), .C1(n132), .C2(n39), .A(n133), .ZN(
        B[13]) );
  NAND2_X1 U17 ( .A1(n104), .A2(n349), .ZN(n74) );
  NOR2_X1 U18 ( .A1(n349), .A2(n141), .ZN(n127) );
  BUF_X1 U19 ( .A(n81), .Z(n168) );
  BUF_X1 U20 ( .A(n81), .Z(n169) );
  INV_X1 U21 ( .A(n141), .ZN(n103) );
  BUF_X1 U22 ( .A(n81), .Z(n170) );
  NOR2_X1 U23 ( .A1(n342), .A2(n343), .ZN(n158) );
  BUF_X1 U24 ( .A(n348), .Z(n343) );
  INV_X1 U25 ( .A(n48), .ZN(n73) );
  INV_X1 U26 ( .A(n38), .ZN(n69) );
  BUF_X1 U27 ( .A(n347), .Z(n345) );
  BUF_X1 U28 ( .A(n348), .Z(n344) );
  BUF_X1 U29 ( .A(n347), .Z(n346) );
  OAI222_X1 U30 ( .A1(n88), .A2(n36), .B1(n168), .B2(n37), .C1(n89), .C2(n35), 
        .ZN(n98) );
  INV_X1 U31 ( .A(n84), .ZN(n89) );
  OAI22_X1 U32 ( .A1(n89), .A2(n36), .B1(n88), .B2(n37), .ZN(n91) );
  AOI222_X1 U33 ( .A1(n59), .A2(n103), .B1(n108), .B2(n104), .C1(n117), .C2(
        n341), .ZN(n75) );
  AOI222_X1 U34 ( .A1(n105), .A2(n104), .B1(n99), .B2(n107), .C1(n53), .C2(
        n103), .ZN(n71) );
  AOI222_X1 U35 ( .A1(n102), .A2(n104), .B1(n98), .B2(n107), .C1(n47), .C2(
        n103), .ZN(n67) );
  AOI222_X1 U36 ( .A1(n109), .A2(n104), .B1(n91), .B2(n107), .C1(n110), .C2(
        n103), .ZN(n61) );
  AOI222_X1 U37 ( .A1(n106), .A2(n104), .B1(n90), .B2(n107), .C1(n108), .C2(
        n103), .ZN(n55) );
  AOI221_X1 U38 ( .B1(n85), .B2(A[8]), .C1(n86), .C2(A[7]), .A(n116), .ZN(n66)
         );
  OAI22_X1 U39 ( .A1(n354), .A2(n88), .B1(n353), .B2(n89), .ZN(n116) );
  AOI221_X1 U40 ( .B1(n85), .B2(A[9]), .C1(n86), .C2(A[8]), .A(n97), .ZN(n60)
         );
  OAI22_X1 U41 ( .A1(n355), .A2(n88), .B1(n354), .B2(n89), .ZN(n97) );
  AOI221_X1 U42 ( .B1(n85), .B2(A[10]), .C1(n86), .C2(A[9]), .A(n87), .ZN(n54)
         );
  OAI22_X1 U43 ( .A1(n356), .A2(n88), .B1(n355), .B2(n89), .ZN(n87) );
  AOI221_X1 U44 ( .B1(n85), .B2(A[11]), .C1(n86), .C2(A[10]), .A(n157), .ZN(
        n48) );
  OAI22_X1 U45 ( .A1(n357), .A2(n88), .B1(n356), .B2(n89), .ZN(n157) );
  AOI221_X1 U46 ( .B1(n85), .B2(A[12]), .C1(n86), .C2(A[11]), .A(n114), .ZN(
        n38) );
  OAI22_X1 U47 ( .A1(n358), .A2(n88), .B1(n357), .B2(n89), .ZN(n114) );
  AOI221_X1 U48 ( .B1(n53), .B2(n104), .C1(n52), .C2(n103), .A(n161), .ZN(n123) );
  INV_X1 U49 ( .A(n162), .ZN(n161) );
  AOI22_X1 U50 ( .A1(n120), .A2(n99), .B1(n107), .B2(n105), .ZN(n162) );
  AOI221_X1 U51 ( .B1(n47), .B2(n104), .C1(n45), .C2(n103), .A(n121), .ZN(n111) );
  INV_X1 U52 ( .A(n122), .ZN(n121) );
  AOI22_X1 U53 ( .A1(n120), .A2(n98), .B1(n107), .B2(n102), .ZN(n122) );
  AOI221_X1 U54 ( .B1(n110), .B2(n104), .C1(n65), .C2(n103), .A(n118), .ZN(n92) );
  INV_X1 U55 ( .A(n119), .ZN(n118) );
  AOI22_X1 U56 ( .A1(n120), .A2(n91), .B1(n107), .B2(n109), .ZN(n119) );
  INV_X1 U57 ( .A(n80), .ZN(n85) );
  AOI222_X1 U58 ( .A1(n42), .A2(n64), .B1(n44), .B2(n65), .C1(n46), .C2(n110), 
        .ZN(n149) );
  AOI222_X1 U59 ( .A1(n46), .A2(n102), .B1(n127), .B2(n98), .C1(n44), .C2(n47), 
        .ZN(n133) );
  AOI222_X1 U60 ( .A1(n42), .A2(n73), .B1(n44), .B2(n51), .C1(n46), .C2(n52), 
        .ZN(n72) );
  AOI222_X1 U61 ( .A1(n42), .A2(n69), .B1(n44), .B2(n43), .C1(n46), .C2(n45), 
        .ZN(n68) );
  AOI222_X1 U62 ( .A1(n42), .A2(n63), .B1(n44), .B2(n64), .C1(n46), .C2(n65), 
        .ZN(n62) );
  AOI222_X1 U63 ( .A1(n42), .A2(n51), .B1(n44), .B2(n52), .C1(n46), .C2(n53), 
        .ZN(n50) );
  AOI222_X1 U64 ( .A1(n42), .A2(n43), .B1(n44), .B2(n45), .C1(n46), .C2(n47), 
        .ZN(n41) );
  AOI222_X1 U65 ( .A1(n42), .A2(n57), .B1(n44), .B2(n58), .C1(n46), .C2(n59), 
        .ZN(n56) );
  AOI222_X1 U66 ( .A1(n46), .A2(n109), .B1(n127), .B2(n91), .C1(n44), .C2(n110), .ZN(n130) );
  AOI222_X1 U67 ( .A1(n46), .A2(n106), .B1(n127), .B2(n90), .C1(n44), .C2(n108), .ZN(n126) );
  OAI221_X1 U68 ( .B1(n54), .B2(n74), .C1(n75), .C2(n349), .A(n76), .ZN(B[3])
         );
  OAI221_X1 U69 ( .B1(n70), .B2(n39), .C1(n71), .C2(n349), .A(n72), .ZN(B[4])
         );
  OAI221_X1 U70 ( .B1(n66), .B2(n39), .C1(n67), .C2(n349), .A(n68), .ZN(B[5])
         );
  OAI221_X1 U71 ( .B1(n54), .B2(n39), .C1(n55), .C2(n349), .A(n56), .ZN(B[7])
         );
  OAI221_X1 U72 ( .B1(n70), .B2(n74), .C1(n123), .C2(n349), .A(n155), .ZN(B[0]) );
  AOI222_X1 U73 ( .A1(n46), .A2(n51), .B1(n77), .B2(n156), .C1(n44), .C2(n73), 
        .ZN(n155) );
  OAI221_X1 U74 ( .B1(n66), .B2(n74), .C1(n111), .C2(n349), .A(n112), .ZN(B[1]) );
  OAI221_X1 U75 ( .B1(n60), .B2(n74), .C1(n92), .C2(n349), .A(n93), .ZN(B[2])
         );
  OAI221_X1 U76 ( .B1(n95), .B2(n39), .C1(n101), .C2(n349), .A(n149), .ZN(
        B[10]) );
  OAI221_X1 U77 ( .B1(n125), .B2(n74), .C1(n79), .C2(n39), .A(n142), .ZN(B[11]) );
  OAI221_X1 U78 ( .B1(n128), .B2(n74), .C1(n129), .C2(n39), .A(n130), .ZN(
        B[14]) );
  OAI221_X1 U79 ( .B1(n124), .B2(n74), .C1(n125), .C2(n39), .A(n126), .ZN(
        B[15]) );
  NOR2_X1 U80 ( .A1(n345), .A2(n123), .ZN(B[16]) );
  NOR2_X1 U81 ( .A1(n345), .A2(n111), .ZN(B[17]) );
  NOR2_X1 U82 ( .A1(n345), .A2(n92), .ZN(B[18]) );
  NOR2_X1 U83 ( .A1(n344), .A2(n75), .ZN(B[19]) );
  NOR2_X1 U84 ( .A1(n346), .A2(n71), .ZN(B[20]) );
  NOR2_X1 U85 ( .A1(n345), .A2(n67), .ZN(B[21]) );
  NOR2_X1 U86 ( .A1(n343), .A2(n61), .ZN(B[22]) );
  NOR2_X1 U87 ( .A1(n344), .A2(n55), .ZN(B[23]) );
  NOR2_X1 U88 ( .A1(n344), .A2(n49), .ZN(B[24]) );
  NOR2_X1 U89 ( .A1(n344), .A2(n40), .ZN(B[25]) );
  NOR2_X1 U90 ( .A1(n343), .A2(n101), .ZN(B[26]) );
  NOR3_X1 U91 ( .A1(n100), .A2(n343), .A3(n341), .ZN(B[27]) );
  AND2_X1 U92 ( .A1(n99), .A2(n77), .ZN(B[28]) );
  AND2_X1 U93 ( .A1(n98), .A2(n77), .ZN(B[29]) );
  AND2_X1 U94 ( .A1(n91), .A2(n77), .ZN(B[30]) );
  AOI221_X1 U95 ( .B1(n46), .B2(n108), .C1(n44), .C2(n59), .A(n143), .ZN(n142)
         );
  NOR3_X1 U96 ( .A1(n349), .A2(n341), .A3(n100), .ZN(n143) );
  AOI221_X1 U97 ( .B1(n52), .B2(n42), .C1(n51), .C2(n77), .A(n139), .ZN(n138)
         );
  INV_X1 U98 ( .A(n140), .ZN(n139) );
  AOI222_X1 U99 ( .A1(n46), .A2(n105), .B1(n127), .B2(n99), .C1(n44), .C2(n53), 
        .ZN(n140) );
  NOR2_X1 U100 ( .A1(n37), .A2(n89), .ZN(n90) );
  AND2_X1 U101 ( .A1(n158), .A2(n340), .ZN(n44) );
  AOI22_X1 U102 ( .A1(n105), .A2(n103), .B1(n99), .B2(n104), .ZN(n49) );
  AOI22_X1 U103 ( .A1(n102), .A2(n103), .B1(n98), .B2(n104), .ZN(n40) );
  AOI22_X1 U104 ( .A1(n109), .A2(n103), .B1(n91), .B2(n104), .ZN(n101) );
  NOR2_X1 U105 ( .A1(n340), .A2(n342), .ZN(n120) );
  INV_X1 U106 ( .A(SH[3]), .ZN(n342) );
  NAND2_X1 U107 ( .A1(SH[1]), .A2(n339), .ZN(n81) );
  NAND2_X1 U108 ( .A1(n340), .A2(n342), .ZN(n141) );
  INV_X1 U109 ( .A(n58), .ZN(n125) );
  INV_X1 U110 ( .A(n95), .ZN(n63) );
  INV_X1 U111 ( .A(n79), .ZN(n57) );
  INV_X1 U112 ( .A(n45), .ZN(n131) );
  INV_X1 U113 ( .A(n59), .ZN(n124) );
  INV_X1 U114 ( .A(n65), .ZN(n128) );
  INV_X1 U115 ( .A(n43), .ZN(n132) );
  INV_X1 U116 ( .A(n64), .ZN(n129) );
  INV_X1 U117 ( .A(n117), .ZN(n100) );
  BUF_X1 U118 ( .A(SH[4]), .Z(n347) );
  BUF_X1 U119 ( .A(SH[4]), .Z(n348) );
  NAND2_X1 U120 ( .A1(SH[1]), .A2(SH[0]), .ZN(n80) );
  OAI221_X1 U121 ( .B1(n80), .B2(n37), .C1(n169), .C2(n36), .A(n164), .ZN(n99)
         );
  AOI22_X1 U122 ( .A1(A[29]), .A2(n83), .B1(A[28]), .B2(n84), .ZN(n164) );
  NOR2_X1 U123 ( .A1(n342), .A2(SH[2]), .ZN(n107) );
  OAI221_X1 U124 ( .B1(n80), .B2(n27), .C1(n169), .C2(n26), .A(n137), .ZN(n45)
         );
  AOI22_X1 U125 ( .A1(A[18]), .A2(n83), .B1(A[17]), .B2(n84), .ZN(n137) );
  OAI221_X1 U126 ( .B1(n80), .B2(n26), .C1(n169), .C2(n25), .A(n165), .ZN(n52)
         );
  AOI22_X1 U127 ( .A1(A[17]), .A2(n83), .B1(A[16]), .B2(n84), .ZN(n165) );
  OAI221_X1 U128 ( .B1(n80), .B2(n23), .C1(n168), .C2(n362), .A(n136), .ZN(n43) );
  AOI22_X1 U129 ( .A1(A[14]), .A2(n83), .B1(A[13]), .B2(n84), .ZN(n136) );
  OAI221_X1 U130 ( .B1(n80), .B2(n24), .C1(n170), .C2(n23), .A(n152), .ZN(n64)
         );
  AOI22_X1 U131 ( .A1(A[15]), .A2(n83), .B1(A[14]), .B2(n84), .ZN(n152) );
  OAI221_X1 U132 ( .B1(n80), .B2(n362), .C1(n168), .C2(n361), .A(n160), .ZN(
        n51) );
  AOI22_X1 U133 ( .A1(A[13]), .A2(n83), .B1(A[12]), .B2(n84), .ZN(n160) );
  OAI221_X1 U134 ( .B1(n80), .B2(n33), .C1(n169), .C2(n32), .A(n163), .ZN(n105) );
  AOI22_X1 U135 ( .A1(A[25]), .A2(n83), .B1(A[24]), .B2(n84), .ZN(n163) );
  OAI221_X1 U136 ( .B1(n80), .B2(n34), .C1(n168), .C2(n33), .A(n135), .ZN(n102) );
  AOI22_X1 U138 ( .A1(A[26]), .A2(n83), .B1(A[25]), .B2(n84), .ZN(n135) );
  OAI221_X1 U139 ( .B1(n80), .B2(n35), .C1(n168), .C2(n34), .A(n153), .ZN(n109) );
  AOI22_X1 U140 ( .A1(A[27]), .A2(n83), .B1(A[26]), .B2(n84), .ZN(n153) );
  OAI221_X1 U141 ( .B1(n80), .B2(n30), .C1(n168), .C2(n29), .A(n134), .ZN(n47)
         );
  INV_X1 U142 ( .A(A[23]), .ZN(n29) );
  AOI22_X1 U143 ( .A1(A[22]), .A2(n83), .B1(A[21]), .B2(n84), .ZN(n134) );
  OAI221_X1 U144 ( .B1(n80), .B2(n31), .C1(n170), .C2(n30), .A(n150), .ZN(n110) );
  AOI22_X1 U145 ( .A1(A[23]), .A2(n83), .B1(A[22]), .B2(n84), .ZN(n150) );
  OAI221_X1 U146 ( .B1(n27), .B2(n88), .C1(n26), .C2(n89), .A(n145), .ZN(n59)
         );
  AOI22_X1 U147 ( .A1(A[22]), .A2(n85), .B1(A[21]), .B2(n86), .ZN(n145) );
  OAI221_X1 U148 ( .B1(n26), .B2(n88), .C1(n25), .C2(n89), .A(n151), .ZN(n65)
         );
  AOI22_X1 U149 ( .A1(A[21]), .A2(n85), .B1(n86), .B2(A[20]), .ZN(n151) );
  OAI221_X1 U150 ( .B1(n88), .B2(n28), .C1(n27), .C2(n89), .A(n166), .ZN(n53)
         );
  INV_X1 U151 ( .A(A[21]), .ZN(n28) );
  AOI22_X1 U152 ( .A1(A[23]), .A2(n85), .B1(A[22]), .B2(n86), .ZN(n166) );
  OAI221_X1 U153 ( .B1(n80), .B2(n32), .C1(n169), .C2(n31), .A(n146), .ZN(n108) );
  AOI22_X1 U154 ( .A1(A[24]), .A2(n83), .B1(A[23]), .B2(n84), .ZN(n146) );
  OAI221_X1 U155 ( .B1(n80), .B2(n25), .C1(n170), .C2(n24), .A(n148), .ZN(n58)
         );
  AOI22_X1 U156 ( .A1(A[16]), .A2(n83), .B1(A[15]), .B2(n84), .ZN(n148) );
  AOI221_X1 U157 ( .B1(n85), .B2(A[7]), .C1(n86), .C2(A[6]), .A(n167), .ZN(n70) );
  OAI22_X1 U158 ( .A1(n353), .A2(n88), .B1(n352), .B2(n89), .ZN(n167) );
  AOI221_X1 U159 ( .B1(n85), .B2(A[13]), .C1(n86), .C2(A[12]), .A(n154), .ZN(
        n95) );
  OAI22_X1 U160 ( .A1(n359), .A2(n88), .B1(n358), .B2(n89), .ZN(n154) );
  AOI221_X1 U161 ( .B1(n85), .B2(A[14]), .C1(n86), .C2(A[13]), .A(n147), .ZN(
        n79) );
  OAI22_X1 U162 ( .A1(n360), .A2(n88), .B1(n359), .B2(n89), .ZN(n147) );
  OAI221_X1 U163 ( .B1(n80), .B2(n36), .C1(n169), .C2(n35), .A(n144), .ZN(n106) );
  AOI22_X1 U164 ( .A1(A[28]), .A2(n83), .B1(A[27]), .B2(n84), .ZN(n144) );
  AOI222_X1 U165 ( .A1(n46), .A2(n43), .B1(n77), .B2(n113), .C1(n44), .C2(n69), 
        .ZN(n112) );
  OAI221_X1 U166 ( .B1(n80), .B2(n352), .C1(n170), .C2(n351), .A(n115), .ZN(
        n113) );
  AOI22_X1 U167 ( .A1(A[2]), .A2(n83), .B1(A[1]), .B2(n84), .ZN(n115) );
  AOI222_X1 U168 ( .A1(n46), .A2(n64), .B1(n77), .B2(n94), .C1(n44), .C2(n63), 
        .ZN(n93) );
  OAI221_X1 U169 ( .B1(n80), .B2(n353), .C1(n170), .C2(n352), .A(n96), .ZN(n94) );
  AOI22_X1 U170 ( .A1(A[3]), .A2(n83), .B1(A[2]), .B2(n84), .ZN(n96) );
  AOI222_X1 U171 ( .A1(n46), .A2(n58), .B1(n77), .B2(n78), .C1(n44), .C2(n57), 
        .ZN(n76) );
  OAI221_X1 U172 ( .B1(n80), .B2(n354), .C1(n170), .C2(n353), .A(n82), .ZN(n78) );
  AOI22_X1 U173 ( .A1(A[4]), .A2(n83), .B1(A[3]), .B2(n84), .ZN(n82) );
  AND2_X1 U174 ( .A1(n77), .A2(n90), .ZN(B[31]) );
  OAI221_X1 U175 ( .B1(n80), .B2(n351), .C1(n168), .C2(n350), .A(n159), .ZN(
        n156) );
  AOI22_X1 U176 ( .A1(A[1]), .A2(n83), .B1(A[0]), .B2(n84), .ZN(n159) );
  AND2_X1 U177 ( .A1(SH[2]), .A2(n158), .ZN(n46) );
  INV_X1 U178 ( .A(A[19]), .ZN(n26) );
  INV_X1 U179 ( .A(A[30]), .ZN(n36) );
  INV_X1 U180 ( .A(A[31]), .ZN(n37) );
  INV_X1 U181 ( .A(A[20]), .ZN(n27) );
  INV_X1 U182 ( .A(A[29]), .ZN(n35) );
  INV_X1 U183 ( .A(A[18]), .ZN(n25) );
  INV_X1 U184 ( .A(A[7]), .ZN(n355) );
  INV_X1 U185 ( .A(A[8]), .ZN(n356) );
  INV_X1 U186 ( .A(A[9]), .ZN(n357) );
  INV_X1 U187 ( .A(A[10]), .ZN(n358) );
  INV_X1 U188 ( .A(A[11]), .ZN(n359) );
  INV_X1 U189 ( .A(A[16]), .ZN(n23) );
  INV_X1 U190 ( .A(A[17]), .ZN(n24) );
  INV_X1 U191 ( .A(A[24]), .ZN(n30) );
  INV_X1 U192 ( .A(A[25]), .ZN(n31) );
  INV_X1 U193 ( .A(A[26]), .ZN(n32) );
  INV_X1 U194 ( .A(A[27]), .ZN(n33) );
  INV_X1 U195 ( .A(A[28]), .ZN(n34) );
  INV_X1 U196 ( .A(SH[0]), .ZN(n339) );
  INV_X1 U197 ( .A(SH[2]), .ZN(n340) );
  INV_X1 U198 ( .A(n342), .ZN(n341) );
  INV_X1 U199 ( .A(A[2]), .ZN(n350) );
  INV_X1 U200 ( .A(A[3]), .ZN(n351) );
  INV_X1 U201 ( .A(A[4]), .ZN(n352) );
  INV_X1 U202 ( .A(A[5]), .ZN(n353) );
  INV_X1 U203 ( .A(A[6]), .ZN(n354) );
  INV_X1 U204 ( .A(A[12]), .ZN(n360) );
  INV_X1 U205 ( .A(A[14]), .ZN(n361) );
  INV_X1 U206 ( .A(A[15]), .ZN(n362) );
endmodule


module SHIFTER_GENERIC_N32_DW_sla_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \A[0] , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383;
  assign B[0] = \A[0] ;
  assign \A[0]  = A[0];

  NOR2_X2 U2 ( .A1(SH[2]), .A2(SH[3]), .ZN(n107) );
  MUX2_X1 U171 ( .A(A[1]), .B(\A[0] ), .S(n68), .Z(n111) );
  NAND2_X1 U3 ( .A1(SH[0]), .A2(n360), .ZN(n67) );
  INV_X1 U4 ( .A(n47), .ZN(n90) );
  INV_X1 U5 ( .A(n368), .ZN(n364) );
  INV_X1 U6 ( .A(n56), .ZN(n70) );
  NAND2_X1 U7 ( .A1(n368), .A2(\A[0] ), .ZN(n39) );
  INV_X1 U8 ( .A(n68), .ZN(n60) );
  OAI21_X1 U9 ( .B1(n367), .B2(n42), .A(n39), .ZN(B[6]) );
  OAI21_X1 U10 ( .B1(n367), .B2(n40), .A(n39), .ZN(B[8]) );
  OAI21_X1 U11 ( .B1(n367), .B2(n38), .A(n39), .ZN(B[9]) );
  OAI21_X1 U12 ( .B1(n366), .B2(n81), .A(n39), .ZN(B[12]) );
  OAI21_X1 U13 ( .B1(n366), .B2(n74), .A(n39), .ZN(B[13]) );
  NAND2_X1 U14 ( .A1(n105), .A2(n364), .ZN(n47) );
  INV_X1 U15 ( .A(n87), .ZN(n52) );
  INV_X1 U16 ( .A(n139), .ZN(n120) );
  BUF_X1 U17 ( .A(n363), .Z(n367) );
  BUF_X1 U18 ( .A(n362), .Z(n365) );
  BUF_X1 U19 ( .A(n362), .Z(n366) );
  BUF_X1 U20 ( .A(n363), .Z(n368) );
  NOR2_X1 U21 ( .A1(n361), .A2(SH[3]), .ZN(n105) );
  INV_X1 U22 ( .A(n57), .ZN(n71) );
  OAI222_X1 U23 ( .A1(n68), .A2(n371), .B1(n370), .B2(n67), .C1(n369), .C2(
        n360), .ZN(n133) );
  NAND2_X1 U24 ( .A1(n107), .A2(n364), .ZN(n87) );
  INV_X1 U25 ( .A(n67), .ZN(n59) );
  AOI221_X1 U26 ( .B1(n111), .B2(n105), .C1(n104), .C2(n107), .A(n120), .ZN(
        n43) );
  AOI221_X1 U27 ( .B1(n133), .B2(n105), .C1(n134), .C2(n107), .A(n120), .ZN(
        n42) );
  AOI221_X1 U28 ( .B1(n126), .B2(n105), .C1(n127), .C2(n107), .A(n120), .ZN(
        n41) );
  AOI221_X1 U29 ( .B1(n118), .B2(n105), .C1(n119), .C2(n107), .A(n120), .ZN(
        n40) );
  AOI221_X1 U30 ( .B1(n104), .B2(n105), .C1(n106), .C2(n107), .A(n108), .ZN(
        n38) );
  INV_X1 U31 ( .A(n109), .ZN(n108) );
  AOI21_X1 U32 ( .B1(n110), .B2(n111), .A(n112), .ZN(n109) );
  AOI221_X1 U33 ( .B1(n134), .B2(n105), .C1(n131), .C2(n107), .A(n179), .ZN(
        n95) );
  INV_X1 U34 ( .A(n180), .ZN(n179) );
  AOI21_X1 U35 ( .B1(n110), .B2(n133), .A(n112), .ZN(n180) );
  AOI221_X1 U36 ( .B1(n127), .B2(n105), .C1(n124), .C2(n107), .A(n174), .ZN(
        n88) );
  INV_X1 U37 ( .A(n175), .ZN(n174) );
  AOI21_X1 U38 ( .B1(n110), .B2(n126), .A(n112), .ZN(n175) );
  AOI221_X1 U39 ( .B1(n119), .B2(n105), .C1(n116), .C2(n107), .A(n169), .ZN(
        n81) );
  INV_X1 U40 ( .A(n170), .ZN(n169) );
  AOI21_X1 U41 ( .B1(n110), .B2(n118), .A(n112), .ZN(n170) );
  AOI221_X1 U42 ( .B1(n106), .B2(n105), .C1(n102), .C2(n107), .A(n164), .ZN(
        n74) );
  INV_X1 U43 ( .A(n165), .ZN(n164) );
  AOI22_X1 U44 ( .A1(n159), .A2(n111), .B1(n110), .B2(n104), .ZN(n165) );
  AOI221_X1 U45 ( .B1(n131), .B2(n105), .C1(n97), .C2(n107), .A(n161), .ZN(n62) );
  INV_X1 U46 ( .A(n162), .ZN(n161) );
  AOI22_X1 U47 ( .A1(n159), .A2(n133), .B1(n110), .B2(n134), .ZN(n162) );
  AOI221_X1 U48 ( .B1(n124), .B2(n105), .C1(n91), .C2(n107), .A(n157), .ZN(n48) );
  INV_X1 U49 ( .A(n158), .ZN(n157) );
  AOI22_X1 U50 ( .A1(n159), .A2(n126), .B1(n110), .B2(n127), .ZN(n158) );
  NAND2_X1 U51 ( .A1(SH[1]), .A2(n359), .ZN(n56) );
  AOI222_X1 U52 ( .A1(n90), .A2(n102), .B1(n54), .B2(n106), .C1(n50), .C2(n104), .ZN(n150) );
  AOI222_X1 U53 ( .A1(n90), .A2(n97), .B1(n54), .B2(n131), .C1(n50), .C2(n134), 
        .ZN(n148) );
  AOI222_X1 U54 ( .A1(n90), .A2(n91), .B1(n54), .B2(n124), .C1(n50), .C2(n127), 
        .ZN(n146) );
  AOI222_X1 U55 ( .A1(n90), .A2(n83), .B1(n54), .B2(n116), .C1(n50), .C2(n119), 
        .ZN(n141) );
  AOI222_X1 U56 ( .A1(n90), .A2(n76), .B1(n54), .B2(n102), .C1(n50), .C2(n106), 
        .ZN(n137) );
  AOI222_X1 U57 ( .A1(n90), .A2(n64), .B1(n54), .B2(n97), .C1(n50), .C2(n131), 
        .ZN(n130) );
  AOI222_X1 U58 ( .A1(n90), .A2(n51), .B1(n54), .B2(n91), .C1(n50), .C2(n124), 
        .ZN(n123) );
  AOI222_X1 U59 ( .A1(n90), .A2(n85), .B1(n54), .B2(n83), .C1(n50), .C2(n116), 
        .ZN(n115) );
  AOI222_X1 U60 ( .A1(n90), .A2(n78), .B1(n54), .B2(n76), .C1(n50), .C2(n102), 
        .ZN(n101) );
  AOI222_X1 U61 ( .A1(n90), .A2(n66), .B1(n54), .B2(n64), .C1(n50), .C2(n97), 
        .ZN(n96) );
  AOI222_X1 U62 ( .A1(n90), .A2(n55), .B1(n54), .B2(n51), .C1(n50), .C2(n91), 
        .ZN(n89) );
  OAI21_X1 U63 ( .B1(n365), .B2(n45), .A(n39), .ZN(B[3]) );
  OAI21_X1 U64 ( .B1(n366), .B2(n44), .A(n39), .ZN(B[4]) );
  OAI21_X1 U65 ( .B1(n367), .B2(n43), .A(n39), .ZN(B[5]) );
  OAI21_X1 U66 ( .B1(n367), .B2(n41), .A(n39), .ZN(B[7]) );
  OAI21_X1 U67 ( .B1(n365), .B2(n145), .A(n39), .ZN(B[1]) );
  OAI21_X1 U68 ( .B1(n365), .B2(n72), .A(n39), .ZN(B[2]) );
  OAI21_X1 U69 ( .B1(n366), .B2(n95), .A(n39), .ZN(B[10]) );
  OAI21_X1 U70 ( .B1(n365), .B2(n88), .A(n39), .ZN(B[11]) );
  OAI21_X1 U71 ( .B1(n365), .B2(n62), .A(n39), .ZN(B[14]) );
  OAI21_X1 U72 ( .B1(n366), .B2(n48), .A(n39), .ZN(B[15]) );
  OAI221_X1 U73 ( .B1(n152), .B2(n47), .C1(n142), .C2(n87), .A(n153), .ZN(
        B[16]) );
  OAI221_X1 U74 ( .B1(n138), .B2(n87), .C1(n145), .C2(n364), .A(n150), .ZN(
        B[17]) );
  OAI221_X1 U75 ( .B1(n132), .B2(n87), .C1(n72), .C2(n364), .A(n148), .ZN(
        B[18]) );
  OAI221_X1 U76 ( .B1(n125), .B2(n87), .C1(n45), .C2(n364), .A(n146), .ZN(
        B[19]) );
  OAI221_X1 U77 ( .B1(n117), .B2(n87), .C1(n44), .C2(n364), .A(n141), .ZN(
        B[20]) );
  OAI221_X1 U78 ( .B1(n103), .B2(n87), .C1(n43), .C2(n364), .A(n137), .ZN(
        B[21]) );
  OAI221_X1 U79 ( .B1(n98), .B2(n87), .C1(n42), .C2(n364), .A(n130), .ZN(B[22]) );
  OAI221_X1 U80 ( .B1(n92), .B2(n87), .C1(n41), .C2(n364), .A(n123), .ZN(B[23]) );
  OAI221_X1 U81 ( .B1(n80), .B2(n87), .C1(n40), .C2(n364), .A(n115), .ZN(B[24]) );
  OAI221_X1 U82 ( .B1(n73), .B2(n87), .C1(n38), .C2(n364), .A(n101), .ZN(B[25]) );
  OAI221_X1 U83 ( .B1(n61), .B2(n87), .C1(n95), .C2(n364), .A(n96), .ZN(B[26])
         );
  OAI221_X1 U84 ( .B1(n46), .B2(n87), .C1(n88), .C2(n364), .A(n89), .ZN(B[27])
         );
  OAI221_X1 U85 ( .B1(n80), .B2(n47), .C1(n81), .C2(n364), .A(n82), .ZN(B[28])
         );
  OAI221_X1 U86 ( .B1(n73), .B2(n47), .C1(n74), .C2(n364), .A(n75), .ZN(B[29])
         );
  OAI221_X1 U87 ( .B1(n61), .B2(n47), .C1(n62), .C2(n364), .A(n63), .ZN(B[30])
         );
  OAI21_X1 U88 ( .B1(n369), .B2(n361), .A(n139), .ZN(n143) );
  AOI221_X1 U89 ( .B1(n50), .B2(n118), .C1(n54), .C2(n119), .A(n154), .ZN(n153) );
  INV_X1 U90 ( .A(n39), .ZN(n154) );
  NOR2_X1 U91 ( .A1(n361), .A2(n139), .ZN(n112) );
  NAND2_X1 U92 ( .A1(n359), .A2(n360), .ZN(n68) );
  AND2_X1 U93 ( .A1(n155), .A2(n361), .ZN(n54) );
  AND2_X1 U94 ( .A1(SH[3]), .A2(n361), .ZN(n110) );
  AOI21_X1 U95 ( .B1(n111), .B2(n107), .A(n143), .ZN(n145) );
  AOI21_X1 U96 ( .B1(n133), .B2(n107), .A(n143), .ZN(n72) );
  AOI21_X1 U97 ( .B1(n126), .B2(n107), .A(n143), .ZN(n45) );
  AOI21_X1 U98 ( .B1(n118), .B2(n107), .A(n143), .ZN(n44) );
  NAND2_X1 U99 ( .A1(SH[3]), .A2(\A[0] ), .ZN(n139) );
  INV_X1 U100 ( .A(n138), .ZN(n76) );
  INV_X1 U101 ( .A(n132), .ZN(n64) );
  INV_X1 U102 ( .A(n125), .ZN(n51) );
  INV_X1 U103 ( .A(n142), .ZN(n83) );
  INV_X1 U104 ( .A(n117), .ZN(n85) );
  INV_X1 U105 ( .A(n103), .ZN(n78) );
  INV_X1 U106 ( .A(n98), .ZN(n66) );
  INV_X1 U107 ( .A(n92), .ZN(n55) );
  INV_X1 U108 ( .A(n116), .ZN(n152) );
  AND2_X1 U109 ( .A1(SH[3]), .A2(n364), .ZN(n155) );
  BUF_X1 U110 ( .A(SH[4]), .Z(n363) );
  BUF_X1 U111 ( .A(SH[4]), .Z(n362) );
  OAI221_X1 U112 ( .B1(n370), .B2(n56), .C1(n369), .C2(n57), .A(n176), .ZN(
        n126) );
  AOI22_X1 U113 ( .A1(n59), .A2(A[2]), .B1(A[3]), .B2(n60), .ZN(n176) );
  OAI221_X1 U114 ( .B1(n67), .B2(n375), .C1(n68), .C2(n376), .A(n173), .ZN(
        n119) );
  AOI22_X1 U115 ( .A1(A[6]), .A2(n70), .B1(A[5]), .B2(n71), .ZN(n173) );
  OAI221_X1 U116 ( .B1(n67), .B2(n372), .C1(n68), .C2(n373), .A(n166), .ZN(
        n104) );
  AOI22_X1 U117 ( .A1(A[3]), .A2(n70), .B1(A[2]), .B2(n71), .ZN(n166) );
  OAI221_X1 U118 ( .B1(n67), .B2(n374), .C1(n68), .C2(n375), .A(n178), .ZN(
        n127) );
  AOI22_X1 U119 ( .A1(A[5]), .A2(n70), .B1(A[4]), .B2(n71), .ZN(n178) );
  OAI221_X1 U120 ( .B1(n67), .B2(n379), .C1(n68), .C2(n380), .A(n172), .ZN(
        n116) );
  AOI22_X1 U121 ( .A1(A[10]), .A2(n70), .B1(A[9]), .B2(n71), .ZN(n172) );
  OAI221_X1 U122 ( .B1(n67), .B2(n376), .C1(n68), .C2(n377), .A(n168), .ZN(
        n106) );
  AOI22_X1 U123 ( .A1(A[7]), .A2(n70), .B1(A[6]), .B2(n71), .ZN(n168) );
  OAI221_X1 U124 ( .B1(n67), .B2(n377), .C1(n68), .C2(n378), .A(n181), .ZN(
        n131) );
  AOI22_X1 U125 ( .A1(A[8]), .A2(n70), .B1(A[7]), .B2(n71), .ZN(n181) );
  OAI221_X1 U126 ( .B1(n67), .B2(n378), .C1(n68), .C2(n379), .A(n177), .ZN(
        n124) );
  AOI22_X1 U127 ( .A1(A[9]), .A2(n70), .B1(A[8]), .B2(n71), .ZN(n177) );
  OAI221_X1 U128 ( .B1(n67), .B2(n380), .C1(n68), .C2(n381), .A(n167), .ZN(
        n102) );
  AOI22_X1 U129 ( .A1(A[11]), .A2(n70), .B1(A[10]), .B2(n71), .ZN(n167) );
  OAI221_X1 U130 ( .B1(n67), .B2(n381), .C1(n68), .C2(n382), .A(n163), .ZN(n97) );
  AOI22_X1 U131 ( .A1(A[12]), .A2(n70), .B1(A[11]), .B2(n71), .ZN(n163) );
  OAI221_X1 U132 ( .B1(n67), .B2(n382), .C1(n68), .C2(n383), .A(n160), .ZN(n91) );
  AOI22_X1 U133 ( .A1(A[13]), .A2(n70), .B1(A[12]), .B2(n71), .ZN(n160) );
  OAI221_X1 U134 ( .B1(n56), .B2(n371), .C1(n370), .C2(n57), .A(n171), .ZN(
        n118) );
  AOI22_X1 U135 ( .A1(n59), .A2(A[3]), .B1(A[4]), .B2(n60), .ZN(n171) );
  AOI221_X1 U136 ( .B1(n59), .B2(A[23]), .C1(n60), .C2(A[24]), .A(n121), .ZN(
        n80) );
  INV_X1 U137 ( .A(n122), .ZN(n121) );
  AOI22_X1 U138 ( .A1(A[22]), .A2(n70), .B1(A[21]), .B2(n71), .ZN(n122) );
  AOI221_X1 U139 ( .B1(n59), .B2(A[24]), .C1(n60), .C2(A[25]), .A(n113), .ZN(
        n73) );
  INV_X1 U140 ( .A(n114), .ZN(n113) );
  AOI22_X1 U141 ( .A1(A[23]), .A2(n70), .B1(A[22]), .B2(n71), .ZN(n114) );
  AOI221_X1 U142 ( .B1(n59), .B2(A[25]), .C1(n60), .C2(A[26]), .A(n99), .ZN(
        n61) );
  INV_X1 U143 ( .A(n100), .ZN(n99) );
  AOI22_X1 U144 ( .A1(A[24]), .A2(n70), .B1(A[23]), .B2(n71), .ZN(n100) );
  AOI221_X1 U145 ( .B1(n59), .B2(A[26]), .C1(n60), .C2(A[27]), .A(n93), .ZN(
        n46) );
  INV_X1 U146 ( .A(n94), .ZN(n93) );
  AOI22_X1 U147 ( .A1(A[25]), .A2(n70), .B1(A[24]), .B2(n71), .ZN(n94) );
  AOI221_X1 U148 ( .B1(n59), .B2(A[16]), .C1(n60), .C2(A[17]), .A(n151), .ZN(
        n138) );
  OAI22_X1 U149 ( .A1(n383), .A2(n56), .B1(n382), .B2(n57), .ZN(n151) );
  AOI221_X1 U150 ( .B1(n59), .B2(A[17]), .C1(n60), .C2(A[18]), .A(n149), .ZN(
        n132) );
  OAI22_X1 U151 ( .A1(n30), .A2(n56), .B1(n383), .B2(n57), .ZN(n149) );
  AOI221_X1 U152 ( .B1(n59), .B2(A[18]), .C1(n60), .C2(A[19]), .A(n147), .ZN(
        n125) );
  OAI22_X1 U153 ( .A1(n31), .A2(n56), .B1(n30), .B2(n57), .ZN(n147) );
  AOI221_X1 U154 ( .B1(n59), .B2(A[19]), .C1(n60), .C2(A[20]), .A(n144), .ZN(
        n117) );
  OAI22_X1 U155 ( .A1(n32), .A2(n56), .B1(n31), .B2(n57), .ZN(n144) );
  AOI221_X1 U156 ( .B1(n59), .B2(A[20]), .C1(n60), .C2(A[21]), .A(n140), .ZN(
        n103) );
  OAI22_X1 U157 ( .A1(n33), .A2(n56), .B1(n32), .B2(n57), .ZN(n140) );
  INV_X1 U158 ( .A(A[19]), .ZN(n33) );
  AOI221_X1 U159 ( .B1(n59), .B2(A[21]), .C1(n60), .C2(A[22]), .A(n135), .ZN(
        n98) );
  INV_X1 U160 ( .A(n136), .ZN(n135) );
  AOI22_X1 U161 ( .A1(A[20]), .A2(n70), .B1(A[19]), .B2(n71), .ZN(n136) );
  AOI221_X1 U162 ( .B1(n59), .B2(A[22]), .C1(n60), .C2(A[23]), .A(n128), .ZN(
        n92) );
  INV_X1 U163 ( .A(n129), .ZN(n128) );
  AOI22_X1 U164 ( .A1(A[21]), .A2(n70), .B1(A[20]), .B2(n71), .ZN(n129) );
  AOI221_X1 U165 ( .B1(n59), .B2(A[15]), .C1(n60), .C2(A[16]), .A(n156), .ZN(
        n142) );
  OAI22_X1 U166 ( .A1(n382), .A2(n56), .B1(n381), .B2(n57), .ZN(n156) );
  NAND2_X1 U167 ( .A1(SH[0]), .A2(SH[1]), .ZN(n57) );
  AOI222_X1 U168 ( .A1(n50), .A2(n83), .B1(n52), .B2(n84), .C1(n54), .C2(n85), 
        .ZN(n82) );
  OAI221_X1 U169 ( .B1(n67), .B2(n34), .C1(n68), .C2(n35), .A(n86), .ZN(n84)
         );
  INV_X1 U170 ( .A(A[27]), .ZN(n34) );
  AOI22_X1 U172 ( .A1(A[26]), .A2(n70), .B1(A[25]), .B2(n71), .ZN(n86) );
  AOI222_X1 U173 ( .A1(n50), .A2(n76), .B1(n52), .B2(n77), .C1(n54), .C2(n78), 
        .ZN(n75) );
  OAI221_X1 U174 ( .B1(n67), .B2(n35), .C1(n68), .C2(n36), .A(n79), .ZN(n77)
         );
  AOI22_X1 U175 ( .A1(A[27]), .A2(n70), .B1(A[26]), .B2(n71), .ZN(n79) );
  AOI222_X1 U176 ( .A1(n50), .A2(n64), .B1(n52), .B2(n65), .C1(n54), .C2(n66), 
        .ZN(n63) );
  OAI221_X1 U177 ( .B1(n67), .B2(n36), .C1(n68), .C2(n37), .A(n69), .ZN(n65)
         );
  INV_X1 U178 ( .A(A[30]), .ZN(n37) );
  AOI22_X1 U179 ( .A1(A[28]), .A2(n70), .B1(A[27]), .B2(n71), .ZN(n69) );
  OAI221_X1 U180 ( .B1(n46), .B2(n47), .C1(n48), .C2(n364), .A(n49), .ZN(B[31]) );
  AOI222_X1 U181 ( .A1(n50), .A2(n51), .B1(n52), .B2(n53), .C1(n54), .C2(n55), 
        .ZN(n49) );
  OAI221_X1 U182 ( .B1(n56), .B2(n36), .C1(n57), .C2(n35), .A(n58), .ZN(n53)
         );
  AOI22_X1 U183 ( .A1(A[30]), .A2(n59), .B1(A[31]), .B2(n60), .ZN(n58) );
  AND2_X1 U184 ( .A1(n155), .A2(SH[2]), .ZN(n50) );
  INV_X1 U185 ( .A(n182), .ZN(n134) );
  AOI221_X1 U186 ( .B1(n70), .B2(A[4]), .C1(A[3]), .C2(n71), .A(n183), .ZN(
        n182) );
  OAI22_X1 U187 ( .A1(n373), .A2(n67), .B1(n374), .B2(n68), .ZN(n183) );
  AND2_X1 U188 ( .A1(SH[2]), .A2(SH[3]), .ZN(n159) );
  INV_X1 U189 ( .A(A[28]), .ZN(n35) );
  INV_X1 U190 ( .A(A[29]), .ZN(n36) );
  INV_X1 U191 ( .A(A[2]), .ZN(n371) );
  INV_X1 U192 ( .A(A[16]), .ZN(n30) );
  INV_X1 U193 ( .A(A[17]), .ZN(n31) );
  INV_X1 U194 ( .A(A[18]), .ZN(n32) );
  INV_X1 U195 ( .A(SH[0]), .ZN(n359) );
  INV_X1 U196 ( .A(SH[1]), .ZN(n360) );
  INV_X1 U197 ( .A(SH[2]), .ZN(n361) );
  INV_X1 U198 ( .A(\A[0] ), .ZN(n369) );
  INV_X1 U199 ( .A(A[1]), .ZN(n370) );
  INV_X1 U200 ( .A(A[4]), .ZN(n372) );
  INV_X1 U201 ( .A(A[5]), .ZN(n373) );
  INV_X1 U202 ( .A(A[6]), .ZN(n374) );
  INV_X1 U203 ( .A(A[7]), .ZN(n375) );
  INV_X1 U204 ( .A(A[8]), .ZN(n376) );
  INV_X1 U205 ( .A(A[9]), .ZN(n377) );
  INV_X1 U206 ( .A(A[10]), .ZN(n378) );
  INV_X1 U207 ( .A(A[11]), .ZN(n379) );
  INV_X1 U208 ( .A(A[12]), .ZN(n380) );
  INV_X1 U209 ( .A(A[13]), .ZN(n381) );
  INV_X1 U210 ( .A(A[14]), .ZN(n382) );
  INV_X1 U211 ( .A(A[15]), .ZN(n383) );
endmodule


module SHIFTER_GENERIC_N32_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] , \ML_int[1][28] ,
         \ML_int[1][27] , \ML_int[1][26] , \ML_int[1][25] , \ML_int[1][24] ,
         \ML_int[1][23] , \ML_int[1][22] , \ML_int[1][21] , \ML_int[1][20] ,
         \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][31] , \ML_int[2][30] , \ML_int[2][29] , \ML_int[2][28] ,
         \ML_int[2][27] , \ML_int[2][26] , \ML_int[2][25] , \ML_int[2][24] ,
         \ML_int[2][23] , \ML_int[2][22] , \ML_int[2][21] , \ML_int[2][20] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][31] , \ML_int[3][30] , \ML_int[3][29] , \ML_int[3][28] ,
         \ML_int[3][27] , \ML_int[3][26] , \ML_int[3][25] , \ML_int[3][24] ,
         \ML_int[3][23] , \ML_int[3][22] , \ML_int[3][21] , \ML_int[3][20] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[3][3] , \ML_int[3][2] , \ML_int[3][1] , \ML_int[3][0] ,
         \ML_int[4][31] , \ML_int[4][30] , \ML_int[4][29] , \ML_int[4][28] ,
         \ML_int[4][27] , \ML_int[4][26] , \ML_int[4][25] , \ML_int[4][24] ,
         \ML_int[4][23] , \ML_int[4][22] , \ML_int[4][21] , \ML_int[4][20] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][16] ,
         \ML_int[4][15] , \ML_int[4][14] , \ML_int[4][13] , \ML_int[4][12] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[4][7] , \ML_int[4][6] , \ML_int[4][5] , \ML_int[4][4] ,
         \ML_int[4][3] , \ML_int[4][2] , \ML_int[4][1] , \ML_int[4][0] , n19,
         n20, n21, n22, n23, n24, n25, n26, n90, n91, n92, n93, n94, n95, n96,
         n97, n98;

  MUX2_X1 M1_4_31 ( .A(\ML_int[4][31] ), .B(\ML_int[4][15] ), .S(n97), .Z(
        B[31]) );
  MUX2_X1 M1_4_30 ( .A(\ML_int[4][30] ), .B(\ML_int[4][14] ), .S(SH[4]), .Z(
        B[30]) );
  MUX2_X1 M1_4_29 ( .A(\ML_int[4][29] ), .B(\ML_int[4][13] ), .S(SH[4]), .Z(
        B[29]) );
  MUX2_X1 M1_4_28 ( .A(\ML_int[4][28] ), .B(\ML_int[4][12] ), .S(SH[4]), .Z(
        B[28]) );
  MUX2_X1 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S(n97), .Z(
        B[27]) );
  MUX2_X1 M1_4_26 ( .A(\ML_int[4][26] ), .B(\ML_int[4][10] ), .S(SH[4]), .Z(
        B[26]) );
  MUX2_X1 M1_4_25 ( .A(\ML_int[4][25] ), .B(\ML_int[4][9] ), .S(n97), .Z(B[25]) );
  MUX2_X1 M1_4_24 ( .A(\ML_int[4][24] ), .B(\ML_int[4][8] ), .S(n97), .Z(B[24]) );
  MUX2_X1 M1_4_23 ( .A(\ML_int[4][23] ), .B(\ML_int[4][7] ), .S(n97), .Z(B[23]) );
  MUX2_X1 M1_4_22 ( .A(\ML_int[4][22] ), .B(\ML_int[4][6] ), .S(n97), .Z(B[22]) );
  MUX2_X1 M1_4_21 ( .A(\ML_int[4][21] ), .B(\ML_int[4][5] ), .S(n97), .Z(B[21]) );
  MUX2_X1 M1_4_20 ( .A(\ML_int[4][20] ), .B(\ML_int[4][4] ), .S(n97), .Z(B[20]) );
  MUX2_X1 M1_4_19 ( .A(\ML_int[4][19] ), .B(\ML_int[4][3] ), .S(SH[4]), .Z(
        B[19]) );
  MUX2_X1 M1_4_18 ( .A(\ML_int[4][18] ), .B(\ML_int[4][2] ), .S(n97), .Z(B[18]) );
  MUX2_X1 M1_4_17 ( .A(\ML_int[4][17] ), .B(\ML_int[4][1] ), .S(SH[4]), .Z(
        B[17]) );
  MUX2_X1 M1_4_16 ( .A(\ML_int[4][16] ), .B(\ML_int[4][0] ), .S(SH[4]), .Z(
        B[16]) );
  MUX2_X1 M1_3_31 ( .A(\ML_int[3][31] ), .B(\ML_int[3][23] ), .S(SH[3]), .Z(
        \ML_int[4][31] ) );
  MUX2_X1 M1_3_30 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S(n95), .Z(
        \ML_int[4][30] ) );
  MUX2_X1 M1_3_29 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S(n95), .Z(
        \ML_int[4][29] ) );
  MUX2_X1 M1_3_28 ( .A(\ML_int[3][28] ), .B(\ML_int[3][20] ), .S(n95), .Z(
        \ML_int[4][28] ) );
  MUX2_X1 M1_3_27 ( .A(\ML_int[3][27] ), .B(\ML_int[3][19] ), .S(SH[3]), .Z(
        \ML_int[4][27] ) );
  MUX2_X1 M1_3_26 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S(n95), .Z(
        \ML_int[4][26] ) );
  MUX2_X1 M1_3_25 ( .A(\ML_int[3][25] ), .B(\ML_int[3][17] ), .S(n95), .Z(
        \ML_int[4][25] ) );
  MUX2_X1 M1_3_24 ( .A(\ML_int[3][24] ), .B(\ML_int[3][16] ), .S(n95), .Z(
        \ML_int[4][24] ) );
  MUX2_X1 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S(n95), .Z(
        \ML_int[4][23] ) );
  MUX2_X1 M1_3_22 ( .A(\ML_int[3][22] ), .B(\ML_int[3][14] ), .S(n95), .Z(
        \ML_int[4][22] ) );
  MUX2_X1 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S(n95), .Z(
        \ML_int[4][21] ) );
  MUX2_X1 M1_3_20 ( .A(\ML_int[3][20] ), .B(\ML_int[3][12] ), .S(n95), .Z(
        \ML_int[4][20] ) );
  MUX2_X1 M1_3_19 ( .A(\ML_int[3][19] ), .B(\ML_int[3][11] ), .S(n95), .Z(
        \ML_int[4][19] ) );
  MUX2_X1 M1_3_18 ( .A(\ML_int[3][18] ), .B(\ML_int[3][10] ), .S(n95), .Z(
        \ML_int[4][18] ) );
  MUX2_X1 M1_3_17 ( .A(\ML_int[3][17] ), .B(\ML_int[3][9] ), .S(n95), .Z(
        \ML_int[4][17] ) );
  MUX2_X1 M1_3_16 ( .A(\ML_int[3][16] ), .B(\ML_int[3][8] ), .S(n95), .Z(
        \ML_int[4][16] ) );
  MUX2_X1 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S(n95), .Z(
        \ML_int[4][15] ) );
  MUX2_X1 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S(n95), .Z(
        \ML_int[4][14] ) );
  MUX2_X1 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S(n95), .Z(
        \ML_int[4][13] ) );
  MUX2_X1 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S(n95), .Z(
        \ML_int[4][12] ) );
  MUX2_X1 M1_3_11 ( .A(\ML_int[3][11] ), .B(\ML_int[3][3] ), .S(n95), .Z(
        \ML_int[4][11] ) );
  MUX2_X1 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S(SH[3]), .Z(
        \ML_int[4][10] ) );
  MUX2_X1 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(SH[3]), .Z(
        \ML_int[4][9] ) );
  MUX2_X1 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S(n95), .Z(
        \ML_int[4][8] ) );
  MUX2_X1 M1_2_31 ( .A(\ML_int[2][31] ), .B(\ML_int[2][27] ), .S(SH[2]), .Z(
        \ML_int[3][31] ) );
  MUX2_X1 M1_2_30 ( .A(\ML_int[2][30] ), .B(\ML_int[2][26] ), .S(SH[2]), .Z(
        \ML_int[3][30] ) );
  MUX2_X1 M1_2_29 ( .A(\ML_int[2][29] ), .B(\ML_int[2][25] ), .S(SH[2]), .Z(
        \ML_int[3][29] ) );
  MUX2_X1 M1_2_28 ( .A(\ML_int[2][28] ), .B(\ML_int[2][24] ), .S(SH[2]), .Z(
        \ML_int[3][28] ) );
  MUX2_X1 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(SH[2]), .Z(
        \ML_int[3][27] ) );
  MUX2_X1 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(SH[2]), .Z(
        \ML_int[3][26] ) );
  MUX2_X1 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(SH[2]), .Z(
        \ML_int[3][25] ) );
  MUX2_X1 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(SH[2]), .Z(
        \ML_int[3][24] ) );
  MUX2_X1 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(SH[2]), .Z(
        \ML_int[3][23] ) );
  MUX2_X1 M1_2_22 ( .A(\ML_int[2][22] ), .B(\ML_int[2][18] ), .S(SH[2]), .Z(
        \ML_int[3][22] ) );
  MUX2_X1 M1_2_21 ( .A(\ML_int[2][21] ), .B(\ML_int[2][17] ), .S(SH[2]), .Z(
        \ML_int[3][21] ) );
  MUX2_X1 M1_2_20 ( .A(\ML_int[2][20] ), .B(\ML_int[2][16] ), .S(SH[2]), .Z(
        \ML_int[3][20] ) );
  MUX2_X1 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S(SH[2]), .Z(
        \ML_int[3][19] ) );
  MUX2_X1 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(SH[2]), .Z(
        \ML_int[3][18] ) );
  MUX2_X1 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(SH[2]), .Z(
        \ML_int[3][17] ) );
  MUX2_X1 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S(SH[2]), .Z(
        \ML_int[3][16] ) );
  MUX2_X1 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S(SH[2]), .Z(
        \ML_int[3][15] ) );
  MUX2_X1 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S(SH[2]), .Z(
        \ML_int[3][14] ) );
  MUX2_X1 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S(SH[2]), .Z(
        \ML_int[3][13] ) );
  MUX2_X1 M1_2_12 ( .A(\ML_int[2][12] ), .B(\ML_int[2][8] ), .S(SH[2]), .Z(
        \ML_int[3][12] ) );
  MUX2_X1 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(SH[2]), .Z(
        \ML_int[3][11] ) );
  MUX2_X1 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(SH[2]), .Z(
        \ML_int[3][10] ) );
  MUX2_X1 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(SH[2]), .Z(
        \ML_int[3][9] ) );
  MUX2_X1 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(SH[2]), .Z(
        \ML_int[3][8] ) );
  MUX2_X1 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(SH[2]), .Z(
        \ML_int[3][7] ) );
  MUX2_X1 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(SH[2]), .Z(
        \ML_int[3][6] ) );
  MUX2_X1 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S(SH[2]), .Z(
        \ML_int[3][5] ) );
  MUX2_X1 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(SH[2]), .Z(
        \ML_int[3][4] ) );
  MUX2_X1 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(n92), .Z(
        \ML_int[2][31] ) );
  MUX2_X1 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S(n91), .Z(
        \ML_int[2][30] ) );
  MUX2_X1 M1_1_29 ( .A(\ML_int[1][29] ), .B(\ML_int[1][27] ), .S(n92), .Z(
        \ML_int[2][29] ) );
  MUX2_X1 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S(n91), .Z(
        \ML_int[2][28] ) );
  MUX2_X1 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S(n92), .Z(
        \ML_int[2][27] ) );
  MUX2_X1 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S(n91), .Z(
        \ML_int[2][26] ) );
  MUX2_X1 M1_1_25 ( .A(\ML_int[1][25] ), .B(\ML_int[1][23] ), .S(n91), .Z(
        \ML_int[2][25] ) );
  MUX2_X1 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(n91), .Z(
        \ML_int[2][24] ) );
  MUX2_X1 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S(n91), .Z(
        \ML_int[2][23] ) );
  MUX2_X1 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(n92), .Z(
        \ML_int[2][22] ) );
  MUX2_X1 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(n91), .Z(
        \ML_int[2][21] ) );
  MUX2_X1 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S(n92), .Z(
        \ML_int[2][20] ) );
  MUX2_X1 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(n91), .Z(
        \ML_int[2][19] ) );
  MUX2_X1 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S(n92), .Z(
        \ML_int[2][18] ) );
  MUX2_X1 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S(n92), .Z(
        \ML_int[2][17] ) );
  MUX2_X1 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(n91), .Z(
        \ML_int[2][16] ) );
  MUX2_X1 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(n92), .Z(
        \ML_int[2][15] ) );
  MUX2_X1 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S(n91), .Z(
        \ML_int[2][14] ) );
  MUX2_X1 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(n91), .Z(
        \ML_int[2][13] ) );
  MUX2_X1 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S(n91), .Z(
        \ML_int[2][12] ) );
  MUX2_X1 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(n91), .Z(
        \ML_int[2][11] ) );
  MUX2_X1 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(n91), .Z(
        \ML_int[2][10] ) );
  MUX2_X1 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(n92), .Z(
        \ML_int[2][9] ) );
  MUX2_X1 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(n92), .Z(
        \ML_int[2][8] ) );
  MUX2_X1 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(n92), .Z(
        \ML_int[2][7] ) );
  MUX2_X1 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(n91), .Z(
        \ML_int[2][6] ) );
  MUX2_X1 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(n92), .Z(
        \ML_int[2][5] ) );
  MUX2_X1 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(n92), .Z(
        \ML_int[2][4] ) );
  MUX2_X1 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(n92), .Z(
        \ML_int[2][3] ) );
  MUX2_X1 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(n92), .Z(
        \ML_int[2][2] ) );
  MUX2_X1 M1_0_31 ( .A(A[31]), .B(A[30]), .S(SH[0]), .Z(\ML_int[1][31] ) );
  MUX2_X1 M1_0_30 ( .A(A[30]), .B(A[29]), .S(SH[0]), .Z(\ML_int[1][30] ) );
  MUX2_X1 M1_0_29 ( .A(A[29]), .B(A[28]), .S(SH[0]), .Z(\ML_int[1][29] ) );
  MUX2_X1 M1_0_28 ( .A(A[28]), .B(A[27]), .S(SH[0]), .Z(\ML_int[1][28] ) );
  MUX2_X1 M1_0_27 ( .A(A[27]), .B(A[26]), .S(SH[0]), .Z(\ML_int[1][27] ) );
  MUX2_X1 M1_0_26 ( .A(A[26]), .B(A[25]), .S(SH[0]), .Z(\ML_int[1][26] ) );
  MUX2_X1 M1_0_25 ( .A(A[25]), .B(A[24]), .S(SH[0]), .Z(\ML_int[1][25] ) );
  MUX2_X1 M1_0_24 ( .A(A[24]), .B(A[23]), .S(SH[0]), .Z(\ML_int[1][24] ) );
  MUX2_X1 M1_0_23 ( .A(A[23]), .B(A[22]), .S(SH[0]), .Z(\ML_int[1][23] ) );
  MUX2_X1 M1_0_22 ( .A(A[22]), .B(A[21]), .S(SH[0]), .Z(\ML_int[1][22] ) );
  MUX2_X1 M1_0_21 ( .A(A[21]), .B(A[20]), .S(SH[0]), .Z(\ML_int[1][21] ) );
  MUX2_X1 M1_0_20 ( .A(A[20]), .B(A[19]), .S(SH[0]), .Z(\ML_int[1][20] ) );
  MUX2_X1 M1_0_19 ( .A(A[19]), .B(A[18]), .S(SH[0]), .Z(\ML_int[1][19] ) );
  MUX2_X1 M1_0_18 ( .A(A[18]), .B(A[17]), .S(SH[0]), .Z(\ML_int[1][18] ) );
  MUX2_X1 M1_0_17 ( .A(A[17]), .B(A[16]), .S(SH[0]), .Z(\ML_int[1][17] ) );
  MUX2_X1 M1_0_16 ( .A(A[16]), .B(A[15]), .S(SH[0]), .Z(\ML_int[1][16] ) );
  MUX2_X1 M1_0_15 ( .A(A[15]), .B(A[14]), .S(SH[0]), .Z(\ML_int[1][15] ) );
  MUX2_X1 M1_0_14 ( .A(A[14]), .B(A[13]), .S(SH[0]), .Z(\ML_int[1][14] ) );
  MUX2_X1 M1_0_13 ( .A(A[13]), .B(A[12]), .S(SH[0]), .Z(\ML_int[1][13] ) );
  MUX2_X1 M1_0_12 ( .A(A[12]), .B(A[11]), .S(SH[0]), .Z(\ML_int[1][12] ) );
  MUX2_X1 M1_0_11 ( .A(A[11]), .B(A[10]), .S(SH[0]), .Z(\ML_int[1][11] ) );
  MUX2_X1 M1_0_10 ( .A(A[10]), .B(A[9]), .S(SH[0]), .Z(\ML_int[1][10] ) );
  MUX2_X1 M1_0_9 ( .A(A[9]), .B(A[8]), .S(SH[0]), .Z(\ML_int[1][9] ) );
  MUX2_X1 M1_0_8 ( .A(A[8]), .B(A[7]), .S(SH[0]), .Z(\ML_int[1][8] ) );
  MUX2_X1 M1_0_7 ( .A(A[7]), .B(A[6]), .S(SH[0]), .Z(\ML_int[1][7] ) );
  MUX2_X1 M1_0_6 ( .A(A[6]), .B(A[5]), .S(SH[0]), .Z(\ML_int[1][6] ) );
  MUX2_X1 M1_0_5 ( .A(A[5]), .B(A[4]), .S(SH[0]), .Z(\ML_int[1][5] ) );
  MUX2_X1 M1_0_4 ( .A(A[4]), .B(A[3]), .S(SH[0]), .Z(\ML_int[1][4] ) );
  MUX2_X1 M1_0_3 ( .A(A[3]), .B(A[2]), .S(SH[0]), .Z(\ML_int[1][3] ) );
  MUX2_X1 M1_0_2 ( .A(A[2]), .B(A[1]), .S(SH[0]), .Z(\ML_int[1][2] ) );
  MUX2_X1 M1_0_1 ( .A(A[1]), .B(A[0]), .S(SH[0]), .Z(\ML_int[1][1] ) );
  INV_X1 U3 ( .A(n26), .ZN(\ML_int[4][0] ) );
  INV_X1 U4 ( .A(n25), .ZN(\ML_int[4][1] ) );
  INV_X1 U5 ( .A(n24), .ZN(\ML_int[4][2] ) );
  INV_X1 U6 ( .A(n23), .ZN(\ML_int[4][3] ) );
  INV_X1 U7 ( .A(n22), .ZN(\ML_int[4][4] ) );
  INV_X1 U8 ( .A(n21), .ZN(\ML_int[4][5] ) );
  INV_X1 U9 ( .A(n20), .ZN(\ML_int[4][6] ) );
  INV_X1 U10 ( .A(n19), .ZN(\ML_int[4][7] ) );
  INV_X1 U11 ( .A(n98), .ZN(n97) );
  NOR2_X1 U12 ( .A1(n97), .A2(n23), .ZN(B[3]) );
  NOR2_X1 U13 ( .A1(n97), .A2(n22), .ZN(B[4]) );
  NOR2_X1 U14 ( .A1(n97), .A2(n21), .ZN(B[5]) );
  NOR2_X1 U15 ( .A1(n97), .A2(n20), .ZN(B[6]) );
  NOR2_X1 U16 ( .A1(n97), .A2(n19), .ZN(B[7]) );
  AND2_X1 U17 ( .A1(\ML_int[4][8] ), .A2(n98), .ZN(B[8]) );
  AND2_X1 U18 ( .A1(\ML_int[4][9] ), .A2(n98), .ZN(B[9]) );
  NOR2_X1 U19 ( .A1(n97), .A2(n26), .ZN(B[0]) );
  NOR2_X1 U20 ( .A1(n97), .A2(n25), .ZN(B[1]) );
  NOR2_X1 U21 ( .A1(n97), .A2(n24), .ZN(B[2]) );
  AND2_X1 U22 ( .A1(\ML_int[4][10] ), .A2(n98), .ZN(B[10]) );
  AND2_X1 U23 ( .A1(\ML_int[4][11] ), .A2(n98), .ZN(B[11]) );
  AND2_X1 U24 ( .A1(\ML_int[4][12] ), .A2(n98), .ZN(B[12]) );
  AND2_X1 U25 ( .A1(\ML_int[4][13] ), .A2(n98), .ZN(B[13]) );
  AND2_X1 U26 ( .A1(\ML_int[4][14] ), .A2(n98), .ZN(B[14]) );
  AND2_X1 U27 ( .A1(\ML_int[4][15] ), .A2(n98), .ZN(B[15]) );
  INV_X1 U28 ( .A(n96), .ZN(n95) );
  INV_X1 U29 ( .A(n93), .ZN(n91) );
  INV_X1 U30 ( .A(n93), .ZN(n92) );
  NAND2_X1 U31 ( .A1(\ML_int[3][0] ), .A2(n96), .ZN(n26) );
  NAND2_X1 U32 ( .A1(\ML_int[3][1] ), .A2(n96), .ZN(n25) );
  NAND2_X1 U33 ( .A1(\ML_int[3][2] ), .A2(n96), .ZN(n24) );
  NAND2_X1 U34 ( .A1(\ML_int[3][3] ), .A2(n96), .ZN(n23) );
  NAND2_X1 U35 ( .A1(\ML_int[3][4] ), .A2(n96), .ZN(n22) );
  NAND2_X1 U36 ( .A1(\ML_int[3][5] ), .A2(n96), .ZN(n21) );
  NAND2_X1 U37 ( .A1(\ML_int[3][6] ), .A2(n96), .ZN(n20) );
  NAND2_X1 U38 ( .A1(\ML_int[3][7] ), .A2(n96), .ZN(n19) );
  INV_X1 U39 ( .A(SH[1]), .ZN(n93) );
  INV_X1 U40 ( .A(SH[4]), .ZN(n98) );
  AND2_X1 U41 ( .A1(\ML_int[2][2] ), .A2(n94), .ZN(\ML_int[3][2] ) );
  AND2_X1 U42 ( .A1(\ML_int[2][3] ), .A2(n94), .ZN(\ML_int[3][3] ) );
  AND2_X1 U43 ( .A1(\ML_int[2][0] ), .A2(n94), .ZN(\ML_int[3][0] ) );
  AND2_X1 U44 ( .A1(\ML_int[2][1] ), .A2(n94), .ZN(\ML_int[3][1] ) );
  AND2_X1 U45 ( .A1(\ML_int[1][0] ), .A2(n93), .ZN(\ML_int[2][0] ) );
  AND2_X1 U46 ( .A1(\ML_int[1][1] ), .A2(n93), .ZN(\ML_int[2][1] ) );
  INV_X1 U47 ( .A(SH[0]), .ZN(n90) );
  INV_X1 U48 ( .A(SH[2]), .ZN(n94) );
  AND2_X1 U49 ( .A1(A[0]), .A2(n90), .ZN(\ML_int[1][0] ) );
  INV_X1 U50 ( .A(SH[3]), .ZN(n96) );
endmodule


module boothmul_N16_M16 ( Am, Bm, Pm );
  input [15:0] Am;
  input [15:0] Bm;
  output [31:0] Pm;
  wire   \negAm[9] , \enc2mux[7][2] , \enc2mux[7][1] , \enc2mux[7][0] ,
         \enc2mux[6][2] , \enc2mux[6][1] , \enc2mux[6][0] , \enc2mux[5][2] ,
         \enc2mux[5][1] , \enc2mux[5][0] , \enc2mux[4][2] , \enc2mux[4][1] ,
         \enc2mux[4][0] , \enc2mux[3][2] , \enc2mux[3][1] , \enc2mux[3][0] ,
         \enc2mux[2][2] , \enc2mux[2][1] , \enc2mux[2][0] , \enc2mux[1][2] ,
         \enc2mux[1][1] , \enc2mux[1][0] , \enc2mux[0][2] , \enc2mux[0][1] ,
         \enc2mux[0][0] , \sig_sum[6][28] , \sig_sum[6][27] , \sig_sum[6][26] ,
         \sig_sum[6][25] , \sig_sum[6][24] , \sig_sum[6][23] ,
         \sig_sum[6][22] , \sig_sum[6][21] , \sig_sum[6][20] ,
         \sig_sum[6][19] , \sig_sum[6][18] , \sig_sum[6][17] ,
         \sig_sum[6][16] , \sig_sum[6][15] , \sig_sum[6][14] ,
         \sig_sum[6][13] , \sig_sum[6][12] , \sig_sum[6][11] ,
         \sig_sum[6][10] , \sig_sum[6][9] , \sig_sum[6][8] , \sig_sum[6][7] ,
         \sig_sum[6][6] , \sig_sum[6][5] , \sig_sum[6][4] , \sig_sum[6][3] ,
         \sig_sum[6][2] , \sig_sum[6][1] , \sig_sum[6][0] , \sig_sum[5][26] ,
         \sig_sum[5][25] , \sig_sum[5][24] , \sig_sum[5][23] ,
         \sig_sum[5][22] , \sig_sum[5][21] , \sig_sum[5][20] ,
         \sig_sum[5][19] , \sig_sum[5][18] , \sig_sum[5][17] ,
         \sig_sum[5][16] , \sig_sum[5][15] , \sig_sum[5][14] ,
         \sig_sum[5][13] , \sig_sum[5][12] , \sig_sum[5][11] ,
         \sig_sum[5][10] , \sig_sum[5][9] , \sig_sum[5][8] , \sig_sum[5][7] ,
         \sig_sum[5][6] , \sig_sum[5][5] , \sig_sum[5][4] , \sig_sum[5][3] ,
         \sig_sum[5][2] , \sig_sum[5][1] , \sig_sum[5][0] , \sig_sum[4][24] ,
         \sig_sum[4][23] , \sig_sum[4][22] , \sig_sum[4][21] ,
         \sig_sum[4][20] , \sig_sum[4][19] , \sig_sum[4][18] ,
         \sig_sum[4][17] , \sig_sum[4][16] , \sig_sum[4][15] ,
         \sig_sum[4][14] , \sig_sum[4][13] , \sig_sum[4][12] ,
         \sig_sum[4][11] , \sig_sum[4][10] , \sig_sum[4][9] , \sig_sum[4][8] ,
         \sig_sum[4][7] , \sig_sum[4][6] , \sig_sum[4][5] , \sig_sum[4][4] ,
         \sig_sum[4][3] , \sig_sum[4][2] , \sig_sum[4][1] , \sig_sum[4][0] ,
         \sig_sum[3][22] , \sig_sum[3][21] , \sig_sum[3][20] ,
         \sig_sum[3][19] , \sig_sum[3][18] , \sig_sum[3][17] ,
         \sig_sum[3][16] , \sig_sum[3][15] , \sig_sum[3][14] ,
         \sig_sum[3][13] , \sig_sum[3][12] , \sig_sum[3][11] ,
         \sig_sum[3][10] , \sig_sum[3][9] , \sig_sum[3][8] , \sig_sum[3][7] ,
         \sig_sum[3][6] , \sig_sum[3][5] , \sig_sum[3][4] , \sig_sum[3][3] ,
         \sig_sum[3][2] , \sig_sum[3][1] , \sig_sum[3][0] , \sig_sum[2][21] ,
         \sig_sum[2][20] , \sig_sum[2][19] , \sig_sum[2][18] ,
         \sig_sum[2][17] , \sig_sum[2][16] , \sig_sum[2][15] ,
         \sig_sum[2][14] , \sig_sum[2][13] , \sig_sum[2][12] ,
         \sig_sum[2][11] , \sig_sum[2][10] , \sig_sum[2][9] , \sig_sum[2][8] ,
         \sig_sum[2][7] , \sig_sum[2][6] , \sig_sum[2][5] , \sig_sum[2][4] ,
         \sig_sum[2][3] , \sig_sum[2][2] , \sig_sum[2][1] , \sig_sum[2][0] ,
         \sig_sum[1][18] , \sig_sum[1][17] , \sig_sum[1][16] ,
         \sig_sum[1][15] , \sig_sum[1][14] , \sig_sum[1][13] ,
         \sig_sum[1][12] , \sig_sum[1][11] , \sig_sum[1][10] , \sig_sum[1][9] ,
         \sig_sum[1][8] , \sig_sum[1][7] , \sig_sum[1][6] , \sig_sum[1][5] ,
         \sig_sum[1][4] , \sig_sum[1][3] , \sig_sum[1][2] , \sig_sum[1][1] ,
         \sig_sum[1][0] , \sig_sum[0][19] , \sig_sum[0][16] , \sig_sum[0][15] ,
         \sig_sum[0][14] , \sig_sum[0][13] , \sig_sum[0][12] ,
         \sig_sum[0][11] , \sig_sum[0][10] , \sig_sum[0][9] , \sig_sum[0][8] ,
         \sig_sum[0][7] , \sig_sum[0][6] , \sig_sum[0][5] , \sig_sum[0][4] ,
         \sig_sum[0][3] , \sig_sum[0][2] , \sig_sum[0][1] , \sig_sum[0][0] ,
         \mux2add[7][31] , \mux2add[7][30] , \mux2add[7][29] ,
         \mux2add[7][28] , \mux2add[7][27] , \mux2add[7][26] ,
         \mux2add[7][25] , \mux2add[7][24] , \mux2add[7][23] ,
         \mux2add[7][22] , \mux2add[7][21] , \mux2add[7][20] ,
         \mux2add[7][19] , \mux2add[7][18] , \mux2add[7][17] ,
         \mux2add[7][16] , \mux2add[7][15] , \mux2add[7][14] ,
         \mux2add[7][13] , \mux2add[7][12] , \mux2add[7][11] ,
         \mux2add[7][10] , \mux2add[7][9] , \mux2add[7][8] , \mux2add[7][7] ,
         \mux2add[7][6] , \mux2add[7][5] , \mux2add[7][4] , \mux2add[7][3] ,
         \mux2add[7][2] , \mux2add[7][1] , \mux2add[7][0] , \mux2add[6][29] ,
         \mux2add[6][28] , \mux2add[6][27] , \mux2add[6][26] ,
         \mux2add[6][25] , \mux2add[6][24] , \mux2add[6][23] ,
         \mux2add[6][22] , \mux2add[6][21] , \mux2add[6][20] ,
         \mux2add[6][19] , \mux2add[6][18] , \mux2add[6][17] ,
         \mux2add[6][16] , \mux2add[6][15] , \mux2add[6][14] ,
         \mux2add[6][13] , \mux2add[6][12] , \mux2add[6][11] ,
         \mux2add[6][10] , \mux2add[6][9] , \mux2add[6][8] , \mux2add[6][7] ,
         \mux2add[6][6] , \mux2add[6][5] , \mux2add[6][4] , \mux2add[6][3] ,
         \mux2add[6][2] , \mux2add[6][1] , \mux2add[6][0] , \mux2add[5][27] ,
         \mux2add[5][26] , \mux2add[5][25] , \mux2add[5][24] ,
         \mux2add[5][23] , \mux2add[5][22] , \mux2add[5][21] ,
         \mux2add[5][20] , \mux2add[5][19] , \mux2add[5][18] ,
         \mux2add[5][17] , \mux2add[5][16] , \mux2add[5][15] ,
         \mux2add[5][14] , \mux2add[5][13] , \mux2add[5][12] ,
         \mux2add[5][11] , \mux2add[5][10] , \mux2add[5][9] , \mux2add[5][8] ,
         \mux2add[5][7] , \mux2add[5][6] , \mux2add[5][5] , \mux2add[5][4] ,
         \mux2add[5][3] , \mux2add[5][2] , \mux2add[5][1] , \mux2add[5][0] ,
         \mux2add[4][25] , \mux2add[4][24] , \mux2add[4][23] ,
         \mux2add[4][22] , \mux2add[4][21] , \mux2add[4][20] ,
         \mux2add[4][19] , \mux2add[4][18] , \mux2add[4][17] ,
         \mux2add[4][16] , \mux2add[4][15] , \mux2add[4][14] ,
         \mux2add[4][13] , \mux2add[4][12] , \mux2add[4][11] ,
         \mux2add[4][10] , \mux2add[4][9] , \mux2add[4][8] , \mux2add[4][7] ,
         \mux2add[4][6] , \mux2add[4][5] , \mux2add[4][4] , \mux2add[4][3] ,
         \mux2add[4][2] , \mux2add[4][1] , \mux2add[4][0] , \mux2add[3][23] ,
         \mux2add[3][22] , \mux2add[3][21] , \mux2add[3][20] ,
         \mux2add[3][19] , \mux2add[3][18] , \mux2add[3][17] ,
         \mux2add[3][16] , \mux2add[3][15] , \mux2add[3][14] ,
         \mux2add[3][13] , \mux2add[3][12] , \mux2add[3][11] ,
         \mux2add[3][10] , \mux2add[3][9] , \mux2add[3][8] , \mux2add[3][7] ,
         \mux2add[3][6] , \mux2add[3][5] , \mux2add[3][4] , \mux2add[3][3] ,
         \mux2add[3][2] , \mux2add[3][1] , \mux2add[3][0] , \mux2add[2][21] ,
         \mux2add[2][20] , \mux2add[2][19] , \mux2add[2][18] ,
         \mux2add[2][17] , \mux2add[2][16] , \mux2add[2][15] ,
         \mux2add[2][14] , \mux2add[2][13] , \mux2add[2][12] ,
         \mux2add[2][11] , \mux2add[2][10] , \mux2add[2][9] , \mux2add[2][8] ,
         \mux2add[2][7] , \mux2add[2][6] , \mux2add[2][5] , \mux2add[2][4] ,
         \mux2add[2][3] , \mux2add[2][2] , \mux2add[2][1] , \mux2add[2][0] ,
         \mux2add[1][19] , \mux2add[1][18] , \mux2add[1][17] ,
         \mux2add[1][16] , \mux2add[1][15] , \mux2add[1][14] ,
         \mux2add[1][13] , \mux2add[1][12] , \mux2add[1][11] ,
         \mux2add[1][10] , \mux2add[1][9] , \mux2add[1][8] , \mux2add[1][7] ,
         \mux2add[1][6] , \mux2add[1][5] , \mux2add[1][4] , \mux2add[1][3] ,
         \mux2add[1][2] , \mux2add[1][1] , \mux2add[1][0] , n4, n5, n9, n12,
         n20, n23, n24, n29, n30, n31, n32, n34, n47, n48, n49, n53, n54, n55,
         n56, n326, n328, n330, n332, n334, n336, n338, n340, n342, n344, n346,
         n348, n350, n352, n354, n356, n362, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405;
  assign n328 = Am[0];
  assign n330 = Am[1];
  assign n332 = Am[2];
  assign n334 = Am[3];
  assign n336 = Am[4];
  assign n338 = Am[5];
  assign n340 = Am[6];
  assign n342 = Am[7];
  assign n344 = Am[8];
  assign n346 = Am[9];
  assign n348 = Am[10];
  assign n350 = Am[11];
  assign n352 = Am[12];
  assign n354 = Am[13];
  assign n356 = Am[14];
  assign n362 = Am[15];

  rcas_N16 sub_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n405, n399, n397, n395, 
        n393, n391, n389, n387, n385, n383, n381, n379, n377, n375, n373, n371}), .add_sub(1'b1), .S({n326, n4, n24, n47, n34, n29, \negAm[9] , n23, n32, n9, 
        n53, n54, n12, n48, n49, n30}) );
  encoder_0 enc_0_1 ( .X({Bm[1:0], 1'b0}), .Y({\enc2mux[0][2] , 
        \enc2mux[0][1] , \enc2mux[0][0] }) );
  mux5to1_N18 mux_0_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n402, 
        n402, n402, n398, n396, n394, n392, n390, n388, n386, n384, n382, n380, 
        n378, n376, n374, n372, n370}), .C({n366, n366, n366, n4, n24, n47, 
        n34, n29, \negAm[9] , n23, n32, n9, n53, n54, n12, n48, n49, n30}), 
        .D({n404, n404, n398, n396, n394, n392, n390, n388, n386, n384, n382, 
        n380, n378, n376, n374, n372, n370, 1'b0}), .E({n368, n368, n4, n24, 
        n47, n34, n29, \negAm[9] , n23, n32, n9, n53, n54, n12, n48, n49, n30, 
        1'b0}), .Y({\sig_sum[0][19] , \sig_sum[0][16] , \sig_sum[0][15] , 
        \sig_sum[0][14] , \sig_sum[0][13] , \sig_sum[0][12] , \sig_sum[0][11] , 
        \sig_sum[0][10] , \sig_sum[0][9] , \sig_sum[0][8] , \sig_sum[0][7] , 
        \sig_sum[0][6] , \sig_sum[0][5] , \sig_sum[0][4] , \sig_sum[0][3] , 
        \sig_sum[0][2] , \sig_sum[0][1] , \sig_sum[0][0] }), .SEL({
        \enc2mux[0][2] , \enc2mux[0][1] , \enc2mux[0][0] }) );
  encoder_7 enc_i_1 ( .X(Bm[3:1]), .Y({\enc2mux[1][2] , \enc2mux[1][1] , 
        \enc2mux[1][0] }) );
  mux5to1_N20 mux_i_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n403, n403, n404, n398, n396, n394, n392, n390, n388, n386, n384, n382, 
        n380, n378, n376, n374, n372, n370, 1'b0, 1'b0}), .C({n367, n366, n366, 
        n4, n24, n47, n34, n29, \negAm[9] , n23, n32, n9, n53, n54, n12, n48, 
        n49, n30, 1'b0, 1'b0}), .D({n403, n403, n398, n396, n394, n392, n390, 
        n388, n386, n384, n382, n380, n378, n376, n374, n372, n370, 1'b0, 1'b0, 
        1'b0}), .E({n366, n366, n4, n24, n47, n34, n29, \negAm[9] , n23, n32, 
        n9, n53, n54, n12, n48, n49, n30, 1'b0, 1'b0, 1'b0}), .Y({
        \mux2add[1][19] , \mux2add[1][18] , \mux2add[1][17] , \mux2add[1][16] , 
        \mux2add[1][15] , \mux2add[1][14] , \mux2add[1][13] , \mux2add[1][12] , 
        \mux2add[1][11] , \mux2add[1][10] , \mux2add[1][9] , \mux2add[1][8] , 
        \mux2add[1][7] , \mux2add[1][6] , \mux2add[1][5] , \mux2add[1][4] , 
        \mux2add[1][3] , \mux2add[1][2] , \mux2add[1][1] , \mux2add[1][0] }), 
        .SEL({\enc2mux[1][2] , \enc2mux[1][1] , \enc2mux[1][0] }) );
  rca_N20 add_i_1 ( .A({\mux2add[1][19] , \mux2add[1][18] , \mux2add[1][17] , 
        \mux2add[1][16] , \mux2add[1][15] , \mux2add[1][14] , \mux2add[1][13] , 
        \mux2add[1][12] , \mux2add[1][11] , \mux2add[1][10] , \mux2add[1][9] , 
        \mux2add[1][8] , \mux2add[1][7] , \mux2add[1][6] , \mux2add[1][5] , 
        \mux2add[1][4] , \mux2add[1][3] , \mux2add[1][2] , \mux2add[1][1] , 
        \mux2add[1][0] }), .B({\sig_sum[0][19] , \sig_sum[0][19] , 
        \sig_sum[0][19] , \sig_sum[0][16] , \sig_sum[0][15] , \sig_sum[0][14] , 
        \sig_sum[0][13] , \sig_sum[0][12] , \sig_sum[0][11] , \sig_sum[0][10] , 
        \sig_sum[0][9] , \sig_sum[0][8] , \sig_sum[0][7] , \sig_sum[0][6] , 
        \sig_sum[0][5] , \sig_sum[0][4] , \sig_sum[0][3] , \sig_sum[0][2] , 
        \sig_sum[0][1] , \sig_sum[0][0] }), .S({n5, \sig_sum[1][18] , 
        \sig_sum[1][17] , \sig_sum[1][16] , \sig_sum[1][15] , \sig_sum[1][14] , 
        \sig_sum[1][13] , \sig_sum[1][12] , \sig_sum[1][11] , \sig_sum[1][10] , 
        \sig_sum[1][9] , \sig_sum[1][8] , \sig_sum[1][7] , \sig_sum[1][6] , 
        \sig_sum[1][5] , \sig_sum[1][4] , \sig_sum[1][3] , \sig_sum[1][2] , 
        \sig_sum[1][1] , \sig_sum[1][0] }) );
  encoder_6 enc_i_2 ( .X(Bm[5:3]), .Y({\enc2mux[2][2] , \enc2mux[2][1] , 
        \enc2mux[2][0] }) );
  mux5to1_N22 mux_i_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({n402, n402, n402, n398, n396, n394, n392, n390, n388, 
        n386, n384, n382, n380, n378, n376, n374, n372, n370, 1'b0, 1'b0, 1'b0, 
        1'b0}), .C({n369, n369, n369, n4, n24, n47, n34, n29, \negAm[9] , n23, 
        n32, n9, n53, n54, n12, n48, n49, n30, 1'b0, 1'b0, 1'b0, 1'b0}), .D({
        n403, n403, n398, n396, n394, n392, n390, n388, n386, n384, n382, n380, 
        n378, n376, n374, n372, n370, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n368, 
        n368, n4, n24, n47, n34, n29, \negAm[9] , n23, n32, n9, n53, n54, n12, 
        n48, n49, n30, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\mux2add[2][21] , 
        \mux2add[2][20] , \mux2add[2][19] , \mux2add[2][18] , \mux2add[2][17] , 
        \mux2add[2][16] , \mux2add[2][15] , \mux2add[2][14] , \mux2add[2][13] , 
        \mux2add[2][12] , \mux2add[2][11] , \mux2add[2][10] , \mux2add[2][9] , 
        \mux2add[2][8] , \mux2add[2][7] , \mux2add[2][6] , \mux2add[2][5] , 
        \mux2add[2][4] , \mux2add[2][3] , \mux2add[2][2] , \mux2add[2][1] , 
        \mux2add[2][0] }), .SEL({\enc2mux[2][2] , \enc2mux[2][1] , 
        \enc2mux[2][0] }) );
  rca_N22 add_i_2 ( .A({\mux2add[2][21] , \mux2add[2][20] , \mux2add[2][19] , 
        \mux2add[2][18] , \mux2add[2][17] , \mux2add[2][16] , \mux2add[2][15] , 
        \mux2add[2][14] , \mux2add[2][13] , \mux2add[2][12] , \mux2add[2][11] , 
        \mux2add[2][10] , \mux2add[2][9] , \mux2add[2][8] , \mux2add[2][7] , 
        \mux2add[2][6] , \mux2add[2][5] , \mux2add[2][4] , \mux2add[2][3] , 
        \mux2add[2][2] , \mux2add[2][1] , \mux2add[2][0] }), .B({n5, n5, n5, 
        \sig_sum[1][18] , \sig_sum[1][17] , \sig_sum[1][16] , \sig_sum[1][15] , 
        \sig_sum[1][14] , \sig_sum[1][13] , \sig_sum[1][12] , \sig_sum[1][11] , 
        \sig_sum[1][10] , \sig_sum[1][9] , \sig_sum[1][8] , \sig_sum[1][7] , 
        \sig_sum[1][6] , \sig_sum[1][5] , \sig_sum[1][4] , \sig_sum[1][3] , 
        \sig_sum[1][2] , \sig_sum[1][1] , \sig_sum[1][0] }), .S({
        \sig_sum[2][21] , \sig_sum[2][20] , \sig_sum[2][19] , \sig_sum[2][18] , 
        \sig_sum[2][17] , \sig_sum[2][16] , \sig_sum[2][15] , \sig_sum[2][14] , 
        \sig_sum[2][13] , \sig_sum[2][12] , \sig_sum[2][11] , \sig_sum[2][10] , 
        \sig_sum[2][9] , \sig_sum[2][8] , \sig_sum[2][7] , \sig_sum[2][6] , 
        \sig_sum[2][5] , \sig_sum[2][4] , \sig_sum[2][3] , \sig_sum[2][2] , 
        \sig_sum[2][1] , \sig_sum[2][0] }) );
  encoder_5 enc_i_3 ( .X(Bm[7:5]), .Y({\enc2mux[3][2] , \enc2mux[3][1] , 
        \enc2mux[3][0] }) );
  mux5to1_N24 mux_i_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .B({n404, n404, n404, n399, n397, n395, n393, 
        n391, n389, n387, n385, n383, n381, n379, n377, n375, n372, n371, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .C({n366, n366, n366, n4, n24, n47, 
        n34, n29, \negAm[9] , n23, n32, n9, n53, n54, n12, n48, n49, n30, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n404, n404, n398, n396, n394, n392, 
        n390, n388, n386, n384, n382, n380, n378, n376, n374, n372, n370, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n366, n366, n4, n24, n47, 
        n34, n29, \negAm[9] , n23, n32, n9, n53, n54, n12, n48, n49, n30, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({\mux2add[3][23] , 
        \mux2add[3][22] , \mux2add[3][21] , \mux2add[3][20] , \mux2add[3][19] , 
        \mux2add[3][18] , \mux2add[3][17] , \mux2add[3][16] , \mux2add[3][15] , 
        \mux2add[3][14] , \mux2add[3][13] , \mux2add[3][12] , \mux2add[3][11] , 
        \mux2add[3][10] , \mux2add[3][9] , \mux2add[3][8] , \mux2add[3][7] , 
        \mux2add[3][6] , \mux2add[3][5] , \mux2add[3][4] , \mux2add[3][3] , 
        \mux2add[3][2] , \mux2add[3][1] , \mux2add[3][0] }), .SEL({
        \enc2mux[3][2] , \enc2mux[3][1] , \enc2mux[3][0] }) );
  rca_N24 add_i_3 ( .A({\mux2add[3][23] , \mux2add[3][22] , \mux2add[3][21] , 
        \mux2add[3][20] , \mux2add[3][19] , \mux2add[3][18] , \mux2add[3][17] , 
        \mux2add[3][16] , \mux2add[3][15] , \mux2add[3][14] , \mux2add[3][13] , 
        \mux2add[3][12] , \mux2add[3][11] , \mux2add[3][10] , \mux2add[3][9] , 
        \mux2add[3][8] , \mux2add[3][7] , \mux2add[3][6] , \mux2add[3][5] , 
        \mux2add[3][4] , \mux2add[3][3] , \mux2add[3][2] , \mux2add[3][1] , 
        \mux2add[3][0] }), .B({\sig_sum[2][21] , \sig_sum[2][21] , 
        \sig_sum[2][21] , \sig_sum[2][20] , \sig_sum[2][19] , \sig_sum[2][18] , 
        \sig_sum[2][17] , \sig_sum[2][16] , \sig_sum[2][15] , \sig_sum[2][14] , 
        \sig_sum[2][13] , \sig_sum[2][12] , \sig_sum[2][11] , \sig_sum[2][10] , 
        \sig_sum[2][9] , \sig_sum[2][8] , \sig_sum[2][7] , \sig_sum[2][6] , 
        \sig_sum[2][5] , \sig_sum[2][4] , \sig_sum[2][3] , \sig_sum[2][2] , 
        \sig_sum[2][1] , \sig_sum[2][0] }), .S({n31, \sig_sum[3][22] , 
        \sig_sum[3][21] , \sig_sum[3][20] , \sig_sum[3][19] , \sig_sum[3][18] , 
        \sig_sum[3][17] , \sig_sum[3][16] , \sig_sum[3][15] , \sig_sum[3][14] , 
        \sig_sum[3][13] , \sig_sum[3][12] , \sig_sum[3][11] , \sig_sum[3][10] , 
        \sig_sum[3][9] , \sig_sum[3][8] , \sig_sum[3][7] , \sig_sum[3][6] , 
        \sig_sum[3][5] , \sig_sum[3][4] , \sig_sum[3][3] , \sig_sum[3][2] , 
        \sig_sum[3][1] , \sig_sum[3][0] }) );
  encoder_4 enc_i_4 ( .X(Bm[9:7]), .Y({\enc2mux[4][2] , \enc2mux[4][1] , 
        \enc2mux[4][0] }) );
  mux5to1_N26 mux_i_4 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n403, n403, n403, n398, n396, 
        n394, n392, n390, n388, n386, n384, n382, n380, n378, n376, n374, n372, 
        n370, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .C({n367, n367, 
        n367, n4, n24, n47, n34, n29, \negAm[9] , n23, n32, n9, n53, n54, n12, 
        n48, n49, n30, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({
        n404, n404, n399, n397, n395, n393, n391, n389, n387, n385, n383, n381, 
        n379, n377, n375, n373, n371, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .E({n368, n368, n4, n24, n47, n34, n29, \negAm[9] , n23, 
        n32, n9, n53, n54, n12, n48, n49, n30, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .Y({\mux2add[4][25] , \mux2add[4][24] , 
        \mux2add[4][23] , \mux2add[4][22] , \mux2add[4][21] , \mux2add[4][20] , 
        \mux2add[4][19] , \mux2add[4][18] , \mux2add[4][17] , \mux2add[4][16] , 
        \mux2add[4][15] , \mux2add[4][14] , \mux2add[4][13] , \mux2add[4][12] , 
        \mux2add[4][11] , \mux2add[4][10] , \mux2add[4][9] , \mux2add[4][8] , 
        \mux2add[4][7] , \mux2add[4][6] , \mux2add[4][5] , \mux2add[4][4] , 
        \mux2add[4][3] , \mux2add[4][2] , \mux2add[4][1] , \mux2add[4][0] }), 
        .SEL({\enc2mux[4][2] , \enc2mux[4][1] , \enc2mux[4][0] }) );
  rca_N26 add_i_4 ( .A({\mux2add[4][25] , \mux2add[4][24] , \mux2add[4][23] , 
        \mux2add[4][22] , \mux2add[4][21] , \mux2add[4][20] , \mux2add[4][19] , 
        \mux2add[4][18] , \mux2add[4][17] , \mux2add[4][16] , \mux2add[4][15] , 
        \mux2add[4][14] , \mux2add[4][13] , \mux2add[4][12] , \mux2add[4][11] , 
        \mux2add[4][10] , \mux2add[4][9] , \mux2add[4][8] , \mux2add[4][7] , 
        \mux2add[4][6] , \mux2add[4][5] , \mux2add[4][4] , \mux2add[4][3] , 
        \mux2add[4][2] , \mux2add[4][1] , \mux2add[4][0] }), .B({n31, n31, n31, 
        \sig_sum[3][22] , \sig_sum[3][21] , \sig_sum[3][20] , \sig_sum[3][19] , 
        \sig_sum[3][18] , \sig_sum[3][17] , \sig_sum[3][16] , \sig_sum[3][15] , 
        \sig_sum[3][14] , \sig_sum[3][13] , \sig_sum[3][12] , \sig_sum[3][11] , 
        \sig_sum[3][10] , \sig_sum[3][9] , \sig_sum[3][8] , \sig_sum[3][7] , 
        \sig_sum[3][6] , \sig_sum[3][5] , \sig_sum[3][4] , \sig_sum[3][3] , 
        \sig_sum[3][2] , \sig_sum[3][1] , \sig_sum[3][0] }), .S({n20, 
        \sig_sum[4][24] , \sig_sum[4][23] , \sig_sum[4][22] , \sig_sum[4][21] , 
        \sig_sum[4][20] , \sig_sum[4][19] , \sig_sum[4][18] , \sig_sum[4][17] , 
        \sig_sum[4][16] , \sig_sum[4][15] , \sig_sum[4][14] , \sig_sum[4][13] , 
        \sig_sum[4][12] , \sig_sum[4][11] , \sig_sum[4][10] , \sig_sum[4][9] , 
        \sig_sum[4][8] , \sig_sum[4][7] , \sig_sum[4][6] , \sig_sum[4][5] , 
        \sig_sum[4][4] , \sig_sum[4][3] , \sig_sum[4][2] , \sig_sum[4][1] , 
        \sig_sum[4][0] }) );
  encoder_3 enc_i_5 ( .X(Bm[11:9]), .Y({\enc2mux[5][2] , \enc2mux[5][1] , 
        \enc2mux[5][0] }) );
  mux5to1_N28 mux_i_5 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n403, n403, n402, 
        n398, n396, n394, n392, n390, n388, n386, n384, n382, n380, n378, n376, 
        n374, n372, n370, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .C({n367, n367, n367, n4, n24, n47, n34, n29, \negAm[9] , n23, 
        n32, n9, n53, n54, n12, n48, n49, n30, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .D({n404, n405, n399, n397, n395, n393, 
        n391, n389, n387, n385, n383, n381, n379, n377, n375, n373, n371, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n368, 
        n368, n4, n24, n47, n34, n29, \negAm[9] , n23, n32, n9, n53, n54, n12, 
        n48, n49, n30, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .Y({\mux2add[5][27] , \mux2add[5][26] , \mux2add[5][25] , 
        \mux2add[5][24] , \mux2add[5][23] , \mux2add[5][22] , \mux2add[5][21] , 
        \mux2add[5][20] , \mux2add[5][19] , \mux2add[5][18] , \mux2add[5][17] , 
        \mux2add[5][16] , \mux2add[5][15] , \mux2add[5][14] , \mux2add[5][13] , 
        \mux2add[5][12] , \mux2add[5][11] , \mux2add[5][10] , \mux2add[5][9] , 
        \mux2add[5][8] , \mux2add[5][7] , \mux2add[5][6] , \mux2add[5][5] , 
        \mux2add[5][4] , \mux2add[5][3] , \mux2add[5][2] , \mux2add[5][1] , 
        \mux2add[5][0] }), .SEL({\enc2mux[5][2] , \enc2mux[5][1] , 
        \enc2mux[5][0] }) );
  rca_N28 add_i_5 ( .A({\mux2add[5][27] , \mux2add[5][26] , \mux2add[5][25] , 
        \mux2add[5][24] , \mux2add[5][23] , \mux2add[5][22] , \mux2add[5][21] , 
        \mux2add[5][20] , \mux2add[5][19] , \mux2add[5][18] , \mux2add[5][17] , 
        \mux2add[5][16] , \mux2add[5][15] , \mux2add[5][14] , \mux2add[5][13] , 
        \mux2add[5][12] , \mux2add[5][11] , \mux2add[5][10] , \mux2add[5][9] , 
        \mux2add[5][8] , \mux2add[5][7] , \mux2add[5][6] , \mux2add[5][5] , 
        \mux2add[5][4] , \mux2add[5][3] , \mux2add[5][2] , \mux2add[5][1] , 
        \mux2add[5][0] }), .B({n20, n20, n20, \sig_sum[4][24] , 
        \sig_sum[4][23] , \sig_sum[4][22] , \sig_sum[4][21] , \sig_sum[4][20] , 
        \sig_sum[4][19] , \sig_sum[4][18] , \sig_sum[4][17] , \sig_sum[4][16] , 
        \sig_sum[4][15] , \sig_sum[4][14] , \sig_sum[4][13] , \sig_sum[4][12] , 
        \sig_sum[4][11] , \sig_sum[4][10] , \sig_sum[4][9] , \sig_sum[4][8] , 
        \sig_sum[4][7] , \sig_sum[4][6] , \sig_sum[4][5] , \sig_sum[4][4] , 
        \sig_sum[4][3] , \sig_sum[4][2] , \sig_sum[4][1] , \sig_sum[4][0] }), 
        .S({n56, \sig_sum[5][26] , \sig_sum[5][25] , \sig_sum[5][24] , 
        \sig_sum[5][23] , \sig_sum[5][22] , \sig_sum[5][21] , \sig_sum[5][20] , 
        \sig_sum[5][19] , \sig_sum[5][18] , \sig_sum[5][17] , \sig_sum[5][16] , 
        \sig_sum[5][15] , \sig_sum[5][14] , \sig_sum[5][13] , \sig_sum[5][12] , 
        \sig_sum[5][11] , \sig_sum[5][10] , \sig_sum[5][9] , \sig_sum[5][8] , 
        \sig_sum[5][7] , \sig_sum[5][6] , \sig_sum[5][5] , \sig_sum[5][4] , 
        \sig_sum[5][3] , \sig_sum[5][2] , \sig_sum[5][1] , \sig_sum[5][0] })
         );
  encoder_2 enc_i_6 ( .X(Bm[13:11]), .Y({\enc2mux[6][2] , \enc2mux[6][1] , 
        \enc2mux[6][0] }) );
  mux5to1_N30 mux_i_6 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n402, 
        n402, n402, n398, n396, n394, n392, n390, n388, n386, n384, n382, n380, 
        n378, n376, n374, n372, n370, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .C({n367, n367, n367, n4, n24, n47, 
        n34, n29, \negAm[9] , n23, n32, n9, n53, n54, n12, n48, n49, n30, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .D({n405, n405, n399, n397, n395, n393, n391, n389, n387, n385, n383, 
        n381, n379, n377, n375, n373, n371, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n368, n368, n4, n24, 
        n47, n34, n29, \negAm[9] , n23, n32, n9, n53, n54, n12, n48, n49, n30, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .Y({\mux2add[6][29] , \mux2add[6][28] , \mux2add[6][27] , 
        \mux2add[6][26] , \mux2add[6][25] , \mux2add[6][24] , \mux2add[6][23] , 
        \mux2add[6][22] , \mux2add[6][21] , \mux2add[6][20] , \mux2add[6][19] , 
        \mux2add[6][18] , \mux2add[6][17] , \mux2add[6][16] , \mux2add[6][15] , 
        \mux2add[6][14] , \mux2add[6][13] , \mux2add[6][12] , \mux2add[6][11] , 
        \mux2add[6][10] , \mux2add[6][9] , \mux2add[6][8] , \mux2add[6][7] , 
        \mux2add[6][6] , \mux2add[6][5] , \mux2add[6][4] , \mux2add[6][3] , 
        \mux2add[6][2] , \mux2add[6][1] , \mux2add[6][0] }), .SEL({
        \enc2mux[6][2] , \enc2mux[6][1] , \enc2mux[6][0] }) );
  rca_N30 add_i_6 ( .A({\mux2add[6][29] , \mux2add[6][28] , \mux2add[6][27] , 
        \mux2add[6][26] , \mux2add[6][25] , \mux2add[6][24] , \mux2add[6][23] , 
        \mux2add[6][22] , \mux2add[6][21] , \mux2add[6][20] , \mux2add[6][19] , 
        \mux2add[6][18] , \mux2add[6][17] , \mux2add[6][16] , \mux2add[6][15] , 
        \mux2add[6][14] , \mux2add[6][13] , \mux2add[6][12] , \mux2add[6][11] , 
        \mux2add[6][10] , \mux2add[6][9] , \mux2add[6][8] , \mux2add[6][7] , 
        \mux2add[6][6] , \mux2add[6][5] , \mux2add[6][4] , \mux2add[6][3] , 
        \mux2add[6][2] , \mux2add[6][1] , \mux2add[6][0] }), .B({n56, n56, n56, 
        \sig_sum[5][26] , \sig_sum[5][25] , \sig_sum[5][24] , \sig_sum[5][23] , 
        \sig_sum[5][22] , \sig_sum[5][21] , \sig_sum[5][20] , \sig_sum[5][19] , 
        \sig_sum[5][18] , \sig_sum[5][17] , \sig_sum[5][16] , \sig_sum[5][15] , 
        \sig_sum[5][14] , \sig_sum[5][13] , \sig_sum[5][12] , \sig_sum[5][11] , 
        \sig_sum[5][10] , \sig_sum[5][9] , \sig_sum[5][8] , \sig_sum[5][7] , 
        \sig_sum[5][6] , \sig_sum[5][5] , \sig_sum[5][4] , \sig_sum[5][3] , 
        \sig_sum[5][2] , \sig_sum[5][1] , \sig_sum[5][0] }), .S({n55, 
        \sig_sum[6][28] , \sig_sum[6][27] , \sig_sum[6][26] , \sig_sum[6][25] , 
        \sig_sum[6][24] , \sig_sum[6][23] , \sig_sum[6][22] , \sig_sum[6][21] , 
        \sig_sum[6][20] , \sig_sum[6][19] , \sig_sum[6][18] , \sig_sum[6][17] , 
        \sig_sum[6][16] , \sig_sum[6][15] , \sig_sum[6][14] , \sig_sum[6][13] , 
        \sig_sum[6][12] , \sig_sum[6][11] , \sig_sum[6][10] , \sig_sum[6][9] , 
        \sig_sum[6][8] , \sig_sum[6][7] , \sig_sum[6][6] , \sig_sum[6][5] , 
        \sig_sum[6][4] , \sig_sum[6][3] , \sig_sum[6][2] , \sig_sum[6][1] , 
        \sig_sum[6][0] }) );
  encoder_1 enc_i_7 ( .X(Bm[15:13]), .Y({\enc2mux[7][2] , \enc2mux[7][1] , 
        \enc2mux[7][0] }) );
  mux5to1_N32 mux_i_7 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n403, n402, n402, n398, n396, n394, n392, n390, n388, n386, n384, n382, 
        n380, n378, n376, n374, n372, n370, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .C({n367, n367, n368, 
        n4, n24, n47, n34, n29, \negAm[9] , n23, n32, n9, n53, n54, n12, n48, 
        n49, n30, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .D({n404, n404, n398, n396, n394, n392, n390, 
        n388, n386, n384, n382, n380, n378, n376, n374, n373, n370, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .E({n368, n368, n4, n24, n47, n34, n29, \negAm[9] , n23, n32, 
        n9, n53, n54, n12, n48, n49, n30, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y({
        \mux2add[7][31] , \mux2add[7][30] , \mux2add[7][29] , \mux2add[7][28] , 
        \mux2add[7][27] , \mux2add[7][26] , \mux2add[7][25] , \mux2add[7][24] , 
        \mux2add[7][23] , \mux2add[7][22] , \mux2add[7][21] , \mux2add[7][20] , 
        \mux2add[7][19] , \mux2add[7][18] , \mux2add[7][17] , \mux2add[7][16] , 
        \mux2add[7][15] , \mux2add[7][14] , \mux2add[7][13] , \mux2add[7][12] , 
        \mux2add[7][11] , \mux2add[7][10] , \mux2add[7][9] , \mux2add[7][8] , 
        \mux2add[7][7] , \mux2add[7][6] , \mux2add[7][5] , \mux2add[7][4] , 
        \mux2add[7][3] , \mux2add[7][2] , \mux2add[7][1] , \mux2add[7][0] }), 
        .SEL({\enc2mux[7][2] , \enc2mux[7][1] , \enc2mux[7][0] }) );
  rca_N32 add_i_7 ( .A({\mux2add[7][31] , \mux2add[7][30] , \mux2add[7][29] , 
        \mux2add[7][28] , \mux2add[7][27] , \mux2add[7][26] , \mux2add[7][25] , 
        \mux2add[7][24] , \mux2add[7][23] , \mux2add[7][22] , \mux2add[7][21] , 
        \mux2add[7][20] , \mux2add[7][19] , \mux2add[7][18] , \mux2add[7][17] , 
        \mux2add[7][16] , \mux2add[7][15] , \mux2add[7][14] , \mux2add[7][13] , 
        \mux2add[7][12] , \mux2add[7][11] , \mux2add[7][10] , \mux2add[7][9] , 
        \mux2add[7][8] , \mux2add[7][7] , \mux2add[7][6] , \mux2add[7][5] , 
        \mux2add[7][4] , \mux2add[7][3] , \mux2add[7][2] , \mux2add[7][1] , 
        \mux2add[7][0] }), .B({n55, n55, n55, \sig_sum[6][28] , 
        \sig_sum[6][27] , \sig_sum[6][26] , \sig_sum[6][25] , \sig_sum[6][24] , 
        \sig_sum[6][23] , \sig_sum[6][22] , \sig_sum[6][21] , \sig_sum[6][20] , 
        \sig_sum[6][19] , \sig_sum[6][18] , \sig_sum[6][17] , \sig_sum[6][16] , 
        \sig_sum[6][15] , \sig_sum[6][14] , \sig_sum[6][13] , \sig_sum[6][12] , 
        \sig_sum[6][11] , \sig_sum[6][10] , \sig_sum[6][9] , \sig_sum[6][8] , 
        \sig_sum[6][7] , \sig_sum[6][6] , \sig_sum[6][5] , \sig_sum[6][4] , 
        \sig_sum[6][3] , \sig_sum[6][2] , \sig_sum[6][1] , \sig_sum[6][0] }), 
        .S(Pm) );
  BUF_X1 U3 ( .A(n365), .Z(n368) );
  BUF_X1 U4 ( .A(n401), .Z(n404) );
  BUF_X1 U5 ( .A(n400), .Z(n402) );
  BUF_X1 U6 ( .A(n364), .Z(n366) );
  BUF_X1 U7 ( .A(n400), .Z(n403) );
  BUF_X1 U8 ( .A(n364), .Z(n367) );
  BUF_X1 U9 ( .A(n401), .Z(n405) );
  BUF_X1 U10 ( .A(n365), .Z(n369) );
  BUF_X1 U11 ( .A(n330), .Z(n372) );
  BUF_X1 U12 ( .A(n354), .Z(n396) );
  BUF_X1 U13 ( .A(n352), .Z(n394) );
  BUF_X1 U14 ( .A(n350), .Z(n392) );
  BUF_X1 U15 ( .A(n348), .Z(n390) );
  BUF_X1 U16 ( .A(n346), .Z(n388) );
  BUF_X1 U17 ( .A(n344), .Z(n386) );
  BUF_X1 U18 ( .A(n342), .Z(n384) );
  BUF_X1 U19 ( .A(n340), .Z(n382) );
  BUF_X1 U20 ( .A(n338), .Z(n380) );
  BUF_X1 U21 ( .A(n334), .Z(n376) );
  BUF_X1 U22 ( .A(n356), .Z(n398) );
  BUF_X1 U23 ( .A(n336), .Z(n378) );
  BUF_X1 U24 ( .A(n332), .Z(n374) );
  BUF_X1 U25 ( .A(n328), .Z(n370) );
  BUF_X1 U26 ( .A(n330), .Z(n373) );
  BUF_X1 U27 ( .A(n356), .Z(n399) );
  BUF_X1 U28 ( .A(n354), .Z(n397) );
  BUF_X1 U29 ( .A(n352), .Z(n395) );
  BUF_X1 U30 ( .A(n350), .Z(n393) );
  BUF_X1 U31 ( .A(n348), .Z(n391) );
  BUF_X1 U32 ( .A(n346), .Z(n389) );
  BUF_X1 U33 ( .A(n344), .Z(n387) );
  BUF_X1 U34 ( .A(n342), .Z(n385) );
  BUF_X1 U35 ( .A(n340), .Z(n383) );
  BUF_X1 U36 ( .A(n338), .Z(n381) );
  BUF_X1 U37 ( .A(n336), .Z(n379) );
  BUF_X1 U38 ( .A(n334), .Z(n377) );
  BUF_X1 U39 ( .A(n332), .Z(n375) );
  BUF_X1 U40 ( .A(n328), .Z(n371) );
  BUF_X1 U41 ( .A(n362), .Z(n400) );
  BUF_X1 U42 ( .A(n326), .Z(n364) );
  BUF_X1 U43 ( .A(n362), .Z(n401) );
  BUF_X1 U44 ( .A(n326), .Z(n365) );
endmodule


module SHIFTER_GENERIC_N32 ( A, B, LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE, 
        OUTPUT );
  input [31:0] A;
  input [4:0] B;
  output [31:0] OUTPUT;
  input LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE;
  wire   N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, N66, N67, N68, N69, N70, N105, N106, N107, N108, N109,
         N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131,
         N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142,
         N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153,
         N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164,
         N165, N166, N167, N168, N202, N203, N204, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230,
         N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241,
         N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252,
         N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263,
         N264, N265, n238, n239, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259;
  assign n238 = B[3];
  assign n239 = B[4];

  SHIFTER_GENERIC_N32_DW01_ash_0 C88 ( .A(A), .DATA_TC(1'b0), .SH({n259, n258, 
        B[2:0]}), .SH_TC(1'b0), .B({N265, N264, N263, N262, N261, N260, N259, 
        N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, 
        N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, 
        N234}) );
  SHIFTER_GENERIC_N32_DW_sla_0 C86 ( .A(A), .SH({n259, n258, B[2:0]}), .SH_TC(
        1'b0), .B({N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, 
        N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, 
        N211, N210, N209, N208, N207, N206, N205, N204, N203, N202}) );
  SHIFTER_GENERIC_N32_DW_rash_0 C50 ( .A(A), .DATA_TC(1'b0), .SH({n259, n258, 
        B[2:0]}), .SH_TC(1'b0), .B({N168, N167, N166, N165, N164, N163, N162, 
        N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, 
        N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, 
        N137}) );
  SHIFTER_GENERIC_N32_DW_sra_0 C48 ( .A(A), .SH({n259, n258, B[2:0]}), .SH_TC(
        1'b0), .B({N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, 
        N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105}) );
  SHIFTER_GENERIC_N32_DW_lbsh_0 C10 ( .A(A), .SH({n259, n258, B[2:0]}), 
        .SH_TC(1'b0), .B({N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, 
        N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, 
        N46, N45, N44, N43, N42, N41, N40, N39}) );
  SHIFTER_GENERIC_N32_DW_rbsh_0 C8 ( .A(A), .SH({n259, n258, B[2:0]}), .SH_TC(
        1'b0), .B({N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7}) );
  BUF_X1 U5 ( .A(n238), .Z(n258) );
  AOI222_X1 U6 ( .A1(N208), .A2(n257), .B1(N111), .B2(n254), .C1(N143), .C2(
        n251), .ZN(n29) );
  AOI222_X1 U7 ( .A1(N210), .A2(n257), .B1(N113), .B2(n254), .C1(N145), .C2(
        n251), .ZN(n25) );
  AOI222_X1 U8 ( .A1(N211), .A2(n257), .B1(N114), .B2(n254), .C1(N146), .C2(
        n251), .ZN(n17) );
  AOI222_X1 U9 ( .A1(N214), .A2(n255), .B1(N117), .B2(n252), .C1(N149), .C2(
        n249), .ZN(n79) );
  AOI222_X1 U10 ( .A1(N215), .A2(n255), .B1(N118), .B2(n252), .C1(N150), .C2(
        n249), .ZN(n77) );
  AOI222_X1 U13 ( .A1(N42), .A2(n248), .B1(N237), .B2(n245), .C1(N10), .C2(
        n242), .ZN(n34) );
  AOI222_X1 U14 ( .A1(N43), .A2(n248), .B1(N238), .B2(n245), .C1(N11), .C2(
        n242), .ZN(n32) );
  AOI222_X1 U15 ( .A1(N44), .A2(n248), .B1(N239), .B2(n245), .C1(N12), .C2(
        n242), .ZN(n30) );
  AOI222_X1 U16 ( .A1(N45), .A2(n248), .B1(N240), .B2(n245), .C1(N13), .C2(
        n242), .ZN(n28) );
  AOI222_X1 U17 ( .A1(N46), .A2(n248), .B1(N241), .B2(n245), .C1(N14), .C2(
        n242), .ZN(n26) );
  AOI222_X1 U18 ( .A1(N47), .A2(n248), .B1(N242), .B2(n245), .C1(N15), .C2(
        n242), .ZN(n24) );
  AOI222_X1 U19 ( .A1(N48), .A2(n248), .B1(N243), .B2(n245), .C1(N16), .C2(
        n242), .ZN(n16) );
  AOI222_X1 U20 ( .A1(N39), .A2(n246), .B1(N234), .B2(n243), .C1(N7), .C2(n240), .ZN(n84) );
  AOI222_X1 U21 ( .A1(N40), .A2(n246), .B1(N235), .B2(n243), .C1(N8), .C2(n240), .ZN(n62) );
  AOI222_X1 U22 ( .A1(N41), .A2(n247), .B1(N236), .B2(n244), .C1(N9), .C2(n241), .ZN(n40) );
  AOI222_X1 U23 ( .A1(N49), .A2(n246), .B1(N244), .B2(n243), .C1(N17), .C2(
        n240), .ZN(n82) );
  AOI222_X1 U24 ( .A1(N50), .A2(n246), .B1(N245), .B2(n243), .C1(N18), .C2(
        n240), .ZN(n80) );
  AOI222_X1 U25 ( .A1(N51), .A2(n246), .B1(N246), .B2(n243), .C1(N19), .C2(
        n240), .ZN(n78) );
  AOI222_X1 U26 ( .A1(N52), .A2(n246), .B1(N247), .B2(n243), .C1(N20), .C2(
        n240), .ZN(n76) );
  AOI222_X1 U27 ( .A1(N53), .A2(n246), .B1(N248), .B2(n243), .C1(N21), .C2(
        n240), .ZN(n74) );
  AOI222_X1 U28 ( .A1(N54), .A2(n246), .B1(N249), .B2(n243), .C1(N22), .C2(
        n240), .ZN(n72) );
  AOI222_X1 U29 ( .A1(N55), .A2(n246), .B1(N250), .B2(n243), .C1(N23), .C2(
        n240), .ZN(n70) );
  AOI222_X1 U30 ( .A1(N56), .A2(n246), .B1(N251), .B2(n243), .C1(N24), .C2(
        n240), .ZN(n68) );
  AOI222_X1 U31 ( .A1(N57), .A2(n246), .B1(N252), .B2(n243), .C1(N25), .C2(
        n240), .ZN(n66) );
  AOI222_X1 U32 ( .A1(N58), .A2(n246), .B1(N253), .B2(n243), .C1(N26), .C2(
        n240), .ZN(n64) );
  AOI222_X1 U33 ( .A1(N59), .A2(n247), .B1(N254), .B2(n244), .C1(N27), .C2(
        n241), .ZN(n60) );
  AOI222_X1 U34 ( .A1(N60), .A2(n247), .B1(N255), .B2(n244), .C1(N28), .C2(
        n241), .ZN(n58) );
  AOI222_X1 U35 ( .A1(N61), .A2(n247), .B1(N256), .B2(n244), .C1(N29), .C2(
        n241), .ZN(n56) );
  AOI222_X1 U36 ( .A1(N62), .A2(n247), .B1(N257), .B2(n244), .C1(N30), .C2(
        n241), .ZN(n54) );
  AOI222_X1 U37 ( .A1(N63), .A2(n247), .B1(N258), .B2(n244), .C1(N31), .C2(
        n241), .ZN(n52) );
  AOI222_X1 U38 ( .A1(N64), .A2(n247), .B1(N259), .B2(n244), .C1(N32), .C2(
        n241), .ZN(n50) );
  AOI222_X1 U39 ( .A1(N65), .A2(n247), .B1(N260), .B2(n244), .C1(N33), .C2(
        n241), .ZN(n48) );
  AOI222_X1 U40 ( .A1(N66), .A2(n247), .B1(N261), .B2(n244), .C1(N34), .C2(
        n241), .ZN(n46) );
  AOI222_X1 U41 ( .A1(N67), .A2(n247), .B1(N262), .B2(n244), .C1(N35), .C2(
        n241), .ZN(n44) );
  AOI222_X1 U42 ( .A1(N68), .A2(n247), .B1(N263), .B2(n244), .C1(N36), .C2(
        n241), .ZN(n42) );
  BUF_X1 U43 ( .A(n22), .Z(n243) );
  BUF_X1 U44 ( .A(n22), .Z(n244) );
  BUF_X1 U45 ( .A(n22), .Z(n245) );
  AOI222_X1 U46 ( .A1(N205), .A2(n257), .B1(N108), .B2(n254), .C1(N140), .C2(
        n251), .ZN(n35) );
  AOI222_X1 U47 ( .A1(N206), .A2(n257), .B1(N109), .B2(n254), .C1(N141), .C2(
        n251), .ZN(n33) );
  AOI222_X1 U48 ( .A1(N207), .A2(n257), .B1(N110), .B2(n254), .C1(N142), .C2(
        n251), .ZN(n31) );
  AOI222_X1 U49 ( .A1(N209), .A2(n257), .B1(N112), .B2(n254), .C1(N144), .C2(
        n251), .ZN(n27) );
  AOI222_X1 U50 ( .A1(N202), .A2(n255), .B1(N105), .B2(n252), .C1(N137), .C2(
        n249), .ZN(n85) );
  AOI222_X1 U51 ( .A1(N203), .A2(n255), .B1(N106), .B2(n252), .C1(N138), .C2(
        n249), .ZN(n63) );
  AOI222_X1 U52 ( .A1(N204), .A2(n256), .B1(N107), .B2(n253), .C1(N139), .C2(
        n250), .ZN(n41) );
  AOI222_X1 U53 ( .A1(N212), .A2(n255), .B1(N115), .B2(n252), .C1(N147), .C2(
        n249), .ZN(n83) );
  AOI222_X1 U54 ( .A1(N213), .A2(n255), .B1(N116), .B2(n252), .C1(N148), .C2(
        n249), .ZN(n81) );
  AOI222_X1 U55 ( .A1(N216), .A2(n255), .B1(N119), .B2(n252), .C1(N151), .C2(
        n249), .ZN(n75) );
  AOI222_X1 U56 ( .A1(N217), .A2(n255), .B1(N120), .B2(n252), .C1(N152), .C2(
        n249), .ZN(n73) );
  AOI222_X1 U57 ( .A1(N218), .A2(n255), .B1(N121), .B2(n252), .C1(N153), .C2(
        n249), .ZN(n71) );
  AOI222_X1 U58 ( .A1(N219), .A2(n255), .B1(N122), .B2(n252), .C1(N154), .C2(
        n249), .ZN(n69) );
  AOI222_X1 U59 ( .A1(N220), .A2(n255), .B1(N123), .B2(n252), .C1(N155), .C2(
        n249), .ZN(n67) );
  AOI222_X1 U60 ( .A1(N221), .A2(n255), .B1(N124), .B2(n252), .C1(N156), .C2(
        n249), .ZN(n65) );
  AOI222_X1 U61 ( .A1(N222), .A2(n256), .B1(N125), .B2(n253), .C1(N157), .C2(
        n250), .ZN(n61) );
  AOI222_X1 U62 ( .A1(N223), .A2(n256), .B1(N126), .B2(n253), .C1(N158), .C2(
        n250), .ZN(n59) );
  AOI222_X1 U63 ( .A1(N224), .A2(n256), .B1(N127), .B2(n253), .C1(N159), .C2(
        n250), .ZN(n57) );
  AOI222_X1 U64 ( .A1(N225), .A2(n256), .B1(N128), .B2(n253), .C1(N160), .C2(
        n250), .ZN(n55) );
  AOI222_X1 U65 ( .A1(N226), .A2(n256), .B1(N129), .B2(n253), .C1(N161), .C2(
        n250), .ZN(n53) );
  AOI222_X1 U66 ( .A1(N227), .A2(n256), .B1(N130), .B2(n253), .C1(N162), .C2(
        n250), .ZN(n51) );
  AOI222_X1 U67 ( .A1(N228), .A2(n256), .B1(N131), .B2(n253), .C1(N163), .C2(
        n250), .ZN(n49) );
  AOI222_X1 U68 ( .A1(N229), .A2(n256), .B1(N132), .B2(n253), .C1(N164), .C2(
        n250), .ZN(n47) );
  AOI222_X1 U69 ( .A1(N230), .A2(n256), .B1(N133), .B2(n253), .C1(N165), .C2(
        n250), .ZN(n45) );
  AOI222_X1 U70 ( .A1(N231), .A2(n256), .B1(N134), .B2(n253), .C1(N166), .C2(
        n250), .ZN(n43) );
  AOI222_X1 U71 ( .A1(N232), .A2(n256), .B1(N135), .B2(n253), .C1(N167), .C2(
        n250), .ZN(n39) );
  NOR3_X1 U72 ( .A1(n87), .A2(n86), .A3(n88), .ZN(n22) );
  AOI222_X1 U73 ( .A1(N70), .A2(n248), .B1(N265), .B2(n245), .C1(N38), .C2(
        n242), .ZN(n36) );
  AOI222_X1 U74 ( .A1(N69), .A2(n247), .B1(N264), .B2(n244), .C1(N37), .C2(
        n241), .ZN(n38) );
  BUF_X1 U75 ( .A(n18), .Z(n255) );
  BUF_X1 U76 ( .A(n18), .Z(n256) );
  BUF_X1 U77 ( .A(n19), .Z(n252) );
  BUF_X1 U78 ( .A(n19), .Z(n253) );
  BUF_X1 U79 ( .A(n20), .Z(n249) );
  BUF_X1 U80 ( .A(n20), .Z(n250) );
  BUF_X1 U81 ( .A(n23), .Z(n240) );
  BUF_X1 U82 ( .A(n23), .Z(n241) );
  BUF_X1 U83 ( .A(n21), .Z(n246) );
  BUF_X1 U84 ( .A(n21), .Z(n247) );
  BUF_X1 U85 ( .A(n19), .Z(n254) );
  BUF_X1 U86 ( .A(n20), .Z(n251) );
  BUF_X1 U87 ( .A(n23), .Z(n242) );
  BUF_X1 U88 ( .A(n18), .Z(n257) );
  BUF_X1 U89 ( .A(n21), .Z(n248) );
  AOI222_X1 U90 ( .A1(N233), .A2(n257), .B1(N136), .B2(n254), .C1(N168), .C2(
        n251), .ZN(n37) );
  NOR3_X1 U91 ( .A1(n86), .A2(LEFT_RIGHT), .A3(n87), .ZN(n20) );
  NOR3_X1 U92 ( .A1(LEFT_RIGHT), .A2(LOGIC_ARITH), .A3(n86), .ZN(n19) );
  NOR3_X1 U93 ( .A1(n86), .A2(LOGIC_ARITH), .A3(n88), .ZN(n18) );
  NOR2_X1 U94 ( .A1(LEFT_RIGHT), .A2(SHIFT_ROTATE), .ZN(n23) );
  NOR2_X1 U95 ( .A1(n88), .A2(SHIFT_ROTATE), .ZN(n21) );
  BUF_X1 U96 ( .A(n239), .Z(n259) );
  INV_X1 U97 ( .A(SHIFT_ROTATE), .ZN(n86) );
  INV_X1 U98 ( .A(LEFT_RIGHT), .ZN(n88) );
  INV_X1 U99 ( .A(LOGIC_ARITH), .ZN(n87) );
  NAND2_X1 U100 ( .A1(n34), .A2(n35), .ZN(OUTPUT[3]) );
  NAND2_X1 U101 ( .A1(n32), .A2(n33), .ZN(OUTPUT[4]) );
  NAND2_X1 U102 ( .A1(n30), .A2(n31), .ZN(OUTPUT[5]) );
  NAND2_X1 U103 ( .A1(n28), .A2(n29), .ZN(OUTPUT[6]) );
  NAND2_X1 U104 ( .A1(n26), .A2(n27), .ZN(OUTPUT[7]) );
  NAND2_X1 U105 ( .A1(n24), .A2(n25), .ZN(OUTPUT[8]) );
  NAND2_X1 U106 ( .A1(n16), .A2(n17), .ZN(OUTPUT[9]) );
  NAND2_X1 U107 ( .A1(n36), .A2(n37), .ZN(OUTPUT[31]) );
  NAND2_X1 U108 ( .A1(n38), .A2(n39), .ZN(OUTPUT[30]) );
  NAND2_X1 U109 ( .A1(n84), .A2(n85), .ZN(OUTPUT[0]) );
  NAND2_X1 U110 ( .A1(n62), .A2(n63), .ZN(OUTPUT[1]) );
  NAND2_X1 U111 ( .A1(n40), .A2(n41), .ZN(OUTPUT[2]) );
  NAND2_X1 U112 ( .A1(n82), .A2(n83), .ZN(OUTPUT[10]) );
  NAND2_X1 U113 ( .A1(n80), .A2(n81), .ZN(OUTPUT[11]) );
  NAND2_X1 U114 ( .A1(n78), .A2(n79), .ZN(OUTPUT[12]) );
  NAND2_X1 U115 ( .A1(n76), .A2(n77), .ZN(OUTPUT[13]) );
  NAND2_X1 U116 ( .A1(n74), .A2(n75), .ZN(OUTPUT[14]) );
  NAND2_X1 U117 ( .A1(n72), .A2(n73), .ZN(OUTPUT[15]) );
  NAND2_X1 U118 ( .A1(n70), .A2(n71), .ZN(OUTPUT[16]) );
  NAND2_X1 U119 ( .A1(n68), .A2(n69), .ZN(OUTPUT[17]) );
  NAND2_X1 U120 ( .A1(n66), .A2(n67), .ZN(OUTPUT[18]) );
  NAND2_X1 U121 ( .A1(n64), .A2(n65), .ZN(OUTPUT[19]) );
  NAND2_X1 U122 ( .A1(n60), .A2(n61), .ZN(OUTPUT[20]) );
  NAND2_X1 U123 ( .A1(n58), .A2(n59), .ZN(OUTPUT[21]) );
  NAND2_X1 U124 ( .A1(n56), .A2(n57), .ZN(OUTPUT[22]) );
  NAND2_X1 U125 ( .A1(n54), .A2(n55), .ZN(OUTPUT[23]) );
  NAND2_X1 U126 ( .A1(n52), .A2(n53), .ZN(OUTPUT[24]) );
  NAND2_X1 U127 ( .A1(n50), .A2(n51), .ZN(OUTPUT[25]) );
  NAND2_X1 U128 ( .A1(n48), .A2(n49), .ZN(OUTPUT[26]) );
  NAND2_X1 U129 ( .A1(n46), .A2(n47), .ZN(OUTPUT[27]) );
  NAND2_X1 U130 ( .A1(n44), .A2(n45), .ZN(OUTPUT[28]) );
  NAND2_X1 U131 ( .A1(n42), .A2(n43), .ZN(OUTPUT[29]) );
endmodule


module comparator ( SUB, Cout, ne, ge, le, ee );
  input [31:0] SUB;
  input Cout;
  output ne, ge, le, ee;
  wire   Cout, n2, n3, n4, n5, n6, n7, n8, n9, n10;
  assign ge = Cout;

  INV_X1 U1 ( .A(ne), .ZN(ee) );
  NOR4_X1 U2 ( .A1(SUB[9]), .A2(SUB[8]), .A3(SUB[7]), .A4(SUB[6]), .ZN(n9) );
  NOR4_X1 U3 ( .A1(SUB[5]), .A2(SUB[4]), .A3(SUB[3]), .A4(SUB[30]), .ZN(n8) );
  NOR4_X1 U4 ( .A1(n10), .A2(SUB[0]), .A3(SUB[11]), .A4(SUB[10]), .ZN(n4) );
  OR4_X1 U5 ( .A1(SUB[13]), .A2(SUB[12]), .A3(SUB[15]), .A4(SUB[14]), .ZN(n10)
         );
  NOR4_X1 U6 ( .A1(SUB[2]), .A2(SUB[29]), .A3(SUB[28]), .A4(SUB[27]), .ZN(n7)
         );
  NOR4_X1 U7 ( .A1(SUB[26]), .A2(SUB[25]), .A3(SUB[24]), .A4(SUB[23]), .ZN(n6)
         );
  NAND4_X1 U8 ( .A1(n2), .A2(n3), .A3(n4), .A4(n5), .ZN(ne) );
  AND4_X1 U9 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .ZN(n5) );
  NOR4_X1 U10 ( .A1(SUB[19]), .A2(SUB[18]), .A3(SUB[17]), .A4(SUB[16]), .ZN(n2) );
  NOR4_X1 U11 ( .A1(SUB[22]), .A2(SUB[21]), .A3(SUB[20]), .A4(SUB[1]), .ZN(n3)
         );
  NAND2_X1 U12 ( .A1(Cout), .A2(ne), .ZN(le) );
endmodule


module P4adder_subtr_N32_M4 ( A, B, Y, SEL, Co );
  input [32:1] A;
  input [32:1] B;
  output [32:1] Y;
  input SEL;
  output Co;
  wire   n22, n23, n24, n25;
  wire   [32:1] xor_B;
  assign n22 = SEL;

  XOR2_X1 U1 ( .A(n23), .B(B[9]), .Z(xor_B[9]) );
  XOR2_X1 U2 ( .A(n23), .B(B[8]), .Z(xor_B[8]) );
  XOR2_X1 U3 ( .A(n23), .B(B[7]), .Z(xor_B[7]) );
  XOR2_X1 U4 ( .A(n23), .B(B[6]), .Z(xor_B[6]) );
  XOR2_X1 U5 ( .A(n23), .B(B[5]), .Z(xor_B[5]) );
  XOR2_X1 U6 ( .A(n23), .B(B[4]), .Z(xor_B[4]) );
  XOR2_X1 U7 ( .A(n23), .B(B[3]), .Z(xor_B[3]) );
  XOR2_X1 U8 ( .A(n23), .B(B[32]), .Z(xor_B[32]) );
  XOR2_X1 U9 ( .A(n23), .B(B[31]), .Z(xor_B[31]) );
  XOR2_X1 U10 ( .A(n23), .B(B[30]), .Z(xor_B[30]) );
  XOR2_X1 U11 ( .A(n23), .B(B[2]), .Z(xor_B[2]) );
  XOR2_X1 U12 ( .A(n23), .B(B[29]), .Z(xor_B[29]) );
  XOR2_X1 U13 ( .A(n24), .B(B[28]), .Z(xor_B[28]) );
  XOR2_X1 U14 ( .A(n24), .B(B[27]), .Z(xor_B[27]) );
  XOR2_X1 U15 ( .A(n24), .B(B[26]), .Z(xor_B[26]) );
  XOR2_X1 U16 ( .A(n24), .B(B[25]), .Z(xor_B[25]) );
  XOR2_X1 U17 ( .A(n24), .B(B[24]), .Z(xor_B[24]) );
  XOR2_X1 U18 ( .A(n24), .B(B[23]), .Z(xor_B[23]) );
  XOR2_X1 U19 ( .A(n24), .B(B[22]), .Z(xor_B[22]) );
  XOR2_X1 U20 ( .A(n24), .B(B[21]), .Z(xor_B[21]) );
  XOR2_X1 U21 ( .A(n24), .B(B[20]), .Z(xor_B[20]) );
  XOR2_X1 U22 ( .A(n24), .B(B[1]), .Z(xor_B[1]) );
  XOR2_X1 U23 ( .A(n24), .B(B[19]), .Z(xor_B[19]) );
  XOR2_X1 U24 ( .A(n24), .B(B[18]), .Z(xor_B[18]) );
  XOR2_X1 U25 ( .A(n25), .B(B[17]), .Z(xor_B[17]) );
  XOR2_X1 U26 ( .A(n25), .B(B[16]), .Z(xor_B[16]) );
  XOR2_X1 U27 ( .A(n25), .B(B[15]), .Z(xor_B[15]) );
  XOR2_X1 U28 ( .A(n25), .B(B[14]), .Z(xor_B[14]) );
  XOR2_X1 U29 ( .A(n25), .B(B[13]), .Z(xor_B[13]) );
  XOR2_X1 U30 ( .A(n25), .B(B[12]), .Z(xor_B[12]) );
  XOR2_X1 U31 ( .A(n25), .B(B[11]), .Z(xor_B[11]) );
  XOR2_X1 U32 ( .A(n25), .B(B[10]), .Z(xor_B[10]) );
  P4adder_N32_M4_1 P4add ( .A(A), .B(xor_B), .Y(Y), .Ci(n25), .Co(Co) );
  BUF_X1 U33 ( .A(n22), .Z(n24) );
  BUF_X1 U34 ( .A(n22), .Z(n23) );
  BUF_X1 U35 ( .A(n22), .Z(n25) );
endmodule


module Logic_Unit_N32 ( R1, R2, S1, S2, S3, S0, Y );
  input [31:0] R1;
  input [31:0] R2;
  output [31:0] Y;
  input S1, S2, S3, S0;
  wire   n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n40, n43, n46, \L3[9] , \L3[8] , \L3[7] , \L3[6] , \L3[5] ,
         \L3[4] , \L3[3] , \L3[31] , \L3[30] , \L3[2] , \L3[29] , \L3[28] ,
         \L3[27] , \L3[26] , \L3[25] , \L3[24] , \L3[23] , \L3[22] , \L3[21] ,
         \L3[20] , \L3[1] , \L3[19] , \L3[18] , \L3[17] , \L3[16] , \L3[15] ,
         \L3[14] , \L3[13] , \L3[12] , \L3[11] , \L3[10] , \L3[0] , \L2[9] ,
         \L2[8] , \L2[7] , \L2[6] , \L2[5] , \L2[4] , \L2[3] , \L2[31] ,
         \L2[30] , \L2[2] , \L2[29] , \L2[28] , \L2[27] , \L2[26] , \L2[25] ,
         \L2[24] , \L2[23] , \L2[22] , \L2[21] , \L2[20] , \L2[1] , \L2[19] ,
         \L2[18] , \L2[17] , \L2[16] , \L2[15] , \L2[14] , \L2[13] , \L2[12] ,
         \L2[11] , \L2[10] , \L2[0] , \L1[9] , \L1[8] , \L1[7] , \L1[6] ,
         \L1[5] , \L1[4] , \L1[3] , \L1[31] , \L1[30] , \L1[2] , \L1[29] ,
         \L1[28] , \L1[27] , \L1[26] , \L1[25] , \L1[24] , \L1[23] , \L1[22] ,
         \L1[21] , \L1[20] , \L1[1] , \L1[19] , \L1[18] , \L1[17] , \L1[16] ,
         \L1[15] , \L1[14] , \L1[13] , \L1[12] , \L1[11] , \L1[10] , \L1[0] ,
         \L0[9] , \L0[8] , \L0[7] , \L0[6] , \L0[5] , \L0[4] , \L0[3] ,
         \L0[31] , \L0[30] , \L0[2] , \L0[29] , \L0[28] , \L0[27] , \L0[26] ,
         \L0[25] , \L0[24] , \L0[23] , \L0[22] , \L0[21] , \L0[20] , \L0[1] ,
         \L0[19] , \L0[18] , \L0[17] , \L0[16] , \L0[15] , \L0[14] , \L0[13] ,
         \L0[12] , \L0[11] , \L0[10] , \L0[0] , n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214;
  wire   [31:0] inv_R2;
  assign n40 = S3;
  assign n43 = S2;
  assign n46 = S1;

  NAND3_0 Nand3_1_0 ( .A(S0), .B(n199), .C(n194), .Y(\L0[0] ) );
  NAND3_127 Nand3_2_0 ( .A(n46), .B(n199), .C(R2[0]), .Y(\L1[0] ) );
  NAND3_126 Nand3_3_0 ( .A(n43), .B(R1[0]), .C(n194), .Y(\L2[0] ) );
  NAND3_125 Nand3_4_0 ( .A(n40), .B(R1[0]), .C(R2[0]), .Y(\L3[0] ) );
  NAND4_0 Nand4_0_0 ( .A(\L0[0] ), .B(\L1[0] ), .C(\L2[0] ), .D(\L3[0] ), .Y(
        Y[0]) );
  NAND3_124 Nand3_1_1 ( .A(S0), .B(n200), .C(n195), .Y(\L0[1] ) );
  NAND3_123 Nand3_2_1 ( .A(n46), .B(n200), .C(R2[1]), .Y(\L1[1] ) );
  NAND3_122 Nand3_3_1 ( .A(n43), .B(R1[1]), .C(n195), .Y(\L2[1] ) );
  NAND3_121 Nand3_4_1 ( .A(n40), .B(R1[1]), .C(R2[1]), .Y(\L3[1] ) );
  NAND4_31 Nand4_0_1 ( .A(\L0[1] ), .B(\L1[1] ), .C(\L2[1] ), .D(\L3[1] ), .Y(
        Y[1]) );
  NAND3_120 Nand3_1_2 ( .A(S0), .B(n201), .C(n196), .Y(\L0[2] ) );
  NAND3_119 Nand3_2_2 ( .A(n46), .B(n201), .C(R2[2]), .Y(\L1[2] ) );
  NAND3_118 Nand3_3_2 ( .A(n43), .B(R1[2]), .C(n196), .Y(\L2[2] ) );
  NAND3_117 Nand3_4_2 ( .A(n40), .B(R1[2]), .C(R2[2]), .Y(\L3[2] ) );
  NAND4_30 Nand4_0_2 ( .A(\L0[2] ), .B(\L1[2] ), .C(\L2[2] ), .D(\L3[2] ), .Y(
        Y[2]) );
  NAND3_116 Nand3_1_3 ( .A(S0), .B(n202), .C(n197), .Y(\L0[3] ) );
  NAND3_115 Nand3_2_3 ( .A(n46), .B(n202), .C(R2[3]), .Y(\L1[3] ) );
  NAND3_114 Nand3_3_3 ( .A(n43), .B(R1[3]), .C(n197), .Y(\L2[3] ) );
  NAND3_113 Nand3_4_3 ( .A(n40), .B(R1[3]), .C(R2[3]), .Y(\L3[3] ) );
  NAND4_29 Nand4_0_3 ( .A(\L0[3] ), .B(\L1[3] ), .C(\L2[3] ), .D(\L3[3] ), .Y(
        Y[3]) );
  NAND3_112 Nand3_1_4 ( .A(S0), .B(n203), .C(n198), .Y(\L0[4] ) );
  NAND3_111 Nand3_2_4 ( .A(n46), .B(n203), .C(R2[4]), .Y(\L1[4] ) );
  NAND3_110 Nand3_3_4 ( .A(n43), .B(R1[4]), .C(n198), .Y(\L2[4] ) );
  NAND3_109 Nand3_4_4 ( .A(n40), .B(R1[4]), .C(R2[4]), .Y(\L3[4] ) );
  NAND4_28 Nand4_0_4 ( .A(\L0[4] ), .B(\L1[4] ), .C(\L2[4] ), .D(\L3[4] ), .Y(
        Y[4]) );
  NAND3_108 Nand3_1_5 ( .A(S0), .B(n204), .C(inv_R2[5]), .Y(\L0[5] ) );
  NAND3_107 Nand3_2_5 ( .A(n46), .B(n204), .C(R2[5]), .Y(\L1[5] ) );
  NAND3_106 Nand3_3_5 ( .A(n43), .B(R1[5]), .C(inv_R2[5]), .Y(\L2[5] ) );
  NAND3_105 Nand3_4_5 ( .A(n40), .B(R1[5]), .C(R2[5]), .Y(\L3[5] ) );
  NAND4_27 Nand4_0_5 ( .A(\L0[5] ), .B(\L1[5] ), .C(\L2[5] ), .D(\L3[5] ), .Y(
        Y[5]) );
  NAND3_104 Nand3_1_6 ( .A(S0), .B(n205), .C(inv_R2[6]), .Y(\L0[6] ) );
  NAND3_103 Nand3_2_6 ( .A(n46), .B(n205), .C(R2[6]), .Y(\L1[6] ) );
  NAND3_102 Nand3_3_6 ( .A(n43), .B(R1[6]), .C(inv_R2[6]), .Y(\L2[6] ) );
  NAND3_101 Nand3_4_6 ( .A(n40), .B(R1[6]), .C(R2[6]), .Y(\L3[6] ) );
  NAND4_26 Nand4_0_6 ( .A(\L0[6] ), .B(\L1[6] ), .C(\L2[6] ), .D(\L3[6] ), .Y(
        Y[6]) );
  NAND3_100 Nand3_1_7 ( .A(S0), .B(n206), .C(inv_R2[7]), .Y(\L0[7] ) );
  NAND3_99 Nand3_2_7 ( .A(n46), .B(n206), .C(R2[7]), .Y(\L1[7] ) );
  NAND3_98 Nand3_3_7 ( .A(n43), .B(R1[7]), .C(inv_R2[7]), .Y(\L2[7] ) );
  NAND3_97 Nand3_4_7 ( .A(n40), .B(R1[7]), .C(R2[7]), .Y(\L3[7] ) );
  NAND4_25 Nand4_0_7 ( .A(\L0[7] ), .B(\L1[7] ), .C(\L2[7] ), .D(\L3[7] ), .Y(
        Y[7]) );
  NAND3_96 Nand3_1_8 ( .A(S0), .B(n207), .C(inv_R2[8]), .Y(\L0[8] ) );
  NAND3_95 Nand3_2_8 ( .A(n46), .B(n207), .C(R2[8]), .Y(\L1[8] ) );
  NAND3_94 Nand3_3_8 ( .A(n43), .B(R1[8]), .C(inv_R2[8]), .Y(\L2[8] ) );
  NAND3_93 Nand3_4_8 ( .A(n40), .B(R1[8]), .C(R2[8]), .Y(\L3[8] ) );
  NAND4_24 Nand4_0_8 ( .A(\L0[8] ), .B(\L1[8] ), .C(\L2[8] ), .D(\L3[8] ), .Y(
        Y[8]) );
  NAND3_92 Nand3_1_9 ( .A(S0), .B(n208), .C(inv_R2[9]), .Y(\L0[9] ) );
  NAND3_91 Nand3_2_9 ( .A(n46), .B(n208), .C(R2[9]), .Y(\L1[9] ) );
  NAND3_90 Nand3_3_9 ( .A(n43), .B(R1[9]), .C(inv_R2[9]), .Y(\L2[9] ) );
  NAND3_89 Nand3_4_9 ( .A(n40), .B(R1[9]), .C(R2[9]), .Y(\L3[9] ) );
  NAND4_23 Nand4_0_9 ( .A(\L0[9] ), .B(\L1[9] ), .C(\L2[9] ), .D(\L3[9] ), .Y(
        Y[9]) );
  NAND3_88 Nand3_1_10 ( .A(S0), .B(n209), .C(inv_R2[10]), .Y(\L0[10] ) );
  NAND3_87 Nand3_2_10 ( .A(n46), .B(n209), .C(R2[10]), .Y(\L1[10] ) );
  NAND3_86 Nand3_3_10 ( .A(n43), .B(R1[10]), .C(inv_R2[10]), .Y(\L2[10] ) );
  NAND3_85 Nand3_4_10 ( .A(n40), .B(R1[10]), .C(R2[10]), .Y(\L3[10] ) );
  NAND4_22 Nand4_0_10 ( .A(\L0[10] ), .B(\L1[10] ), .C(\L2[10] ), .D(\L3[10] ), 
        .Y(Y[10]) );
  NAND3_84 Nand3_1_11 ( .A(S0), .B(n210), .C(inv_R2[11]), .Y(\L0[11] ) );
  NAND3_83 Nand3_2_11 ( .A(n46), .B(n210), .C(R2[11]), .Y(\L1[11] ) );
  NAND3_82 Nand3_3_11 ( .A(n43), .B(R1[11]), .C(inv_R2[11]), .Y(\L2[11] ) );
  NAND3_81 Nand3_4_11 ( .A(n40), .B(R1[11]), .C(R2[11]), .Y(\L3[11] ) );
  NAND4_21 Nand4_0_11 ( .A(\L0[11] ), .B(\L1[11] ), .C(\L2[11] ), .D(\L3[11] ), 
        .Y(Y[11]) );
  NAND3_80 Nand3_1_12 ( .A(S0), .B(n211), .C(inv_R2[12]), .Y(\L0[12] ) );
  NAND3_79 Nand3_2_12 ( .A(n46), .B(n211), .C(R2[12]), .Y(\L1[12] ) );
  NAND3_78 Nand3_3_12 ( .A(n43), .B(R1[12]), .C(inv_R2[12]), .Y(\L2[12] ) );
  NAND3_77 Nand3_4_12 ( .A(n40), .B(R1[12]), .C(R2[12]), .Y(\L3[12] ) );
  NAND4_20 Nand4_0_12 ( .A(\L0[12] ), .B(\L1[12] ), .C(\L2[12] ), .D(\L3[12] ), 
        .Y(Y[12]) );
  NAND3_76 Nand3_1_13 ( .A(S0), .B(n212), .C(inv_R2[13]), .Y(\L0[13] ) );
  NAND3_75 Nand3_2_13 ( .A(n46), .B(n212), .C(R2[13]), .Y(\L1[13] ) );
  NAND3_74 Nand3_3_13 ( .A(n43), .B(R1[13]), .C(inv_R2[13]), .Y(\L2[13] ) );
  NAND3_73 Nand3_4_13 ( .A(n40), .B(R1[13]), .C(R2[13]), .Y(\L3[13] ) );
  NAND4_19 Nand4_0_13 ( .A(\L0[13] ), .B(\L1[13] ), .C(\L2[13] ), .D(\L3[13] ), 
        .Y(Y[13]) );
  NAND3_72 Nand3_1_14 ( .A(S0), .B(n213), .C(inv_R2[14]), .Y(\L0[14] ) );
  NAND3_71 Nand3_2_14 ( .A(n46), .B(n213), .C(R2[14]), .Y(\L1[14] ) );
  NAND3_70 Nand3_3_14 ( .A(n43), .B(R1[14]), .C(inv_R2[14]), .Y(\L2[14] ) );
  NAND3_69 Nand3_4_14 ( .A(n40), .B(R1[14]), .C(R2[14]), .Y(\L3[14] ) );
  NAND4_18 Nand4_0_14 ( .A(\L0[14] ), .B(\L1[14] ), .C(\L2[14] ), .D(\L3[14] ), 
        .Y(Y[14]) );
  NAND3_68 Nand3_1_15 ( .A(S0), .B(n214), .C(inv_R2[15]), .Y(\L0[15] ) );
  NAND3_67 Nand3_2_15 ( .A(n46), .B(n214), .C(R2[15]), .Y(\L1[15] ) );
  NAND3_66 Nand3_3_15 ( .A(n43), .B(R1[15]), .C(inv_R2[15]), .Y(\L2[15] ) );
  NAND3_65 Nand3_4_15 ( .A(n40), .B(R1[15]), .C(R2[15]), .Y(\L3[15] ) );
  NAND4_17 Nand4_0_15 ( .A(\L0[15] ), .B(\L1[15] ), .C(\L2[15] ), .D(\L3[15] ), 
        .Y(Y[15]) );
  NAND3_64 Nand3_1_16 ( .A(S0), .B(n22), .C(inv_R2[16]), .Y(\L0[16] ) );
  NAND3_63 Nand3_2_16 ( .A(n46), .B(n22), .C(R2[16]), .Y(\L1[16] ) );
  NAND3_62 Nand3_3_16 ( .A(n43), .B(R1[16]), .C(inv_R2[16]), .Y(\L2[16] ) );
  NAND3_61 Nand3_4_16 ( .A(n40), .B(R1[16]), .C(R2[16]), .Y(\L3[16] ) );
  NAND4_16 Nand4_0_16 ( .A(\L0[16] ), .B(\L1[16] ), .C(\L2[16] ), .D(\L3[16] ), 
        .Y(Y[16]) );
  NAND3_60 Nand3_1_17 ( .A(S0), .B(n23), .C(inv_R2[17]), .Y(\L0[17] ) );
  NAND3_59 Nand3_2_17 ( .A(n46), .B(n23), .C(R2[17]), .Y(\L1[17] ) );
  NAND3_58 Nand3_3_17 ( .A(n43), .B(R1[17]), .C(inv_R2[17]), .Y(\L2[17] ) );
  NAND3_57 Nand3_4_17 ( .A(n40), .B(R1[17]), .C(R2[17]), .Y(\L3[17] ) );
  NAND4_15 Nand4_0_17 ( .A(\L0[17] ), .B(\L1[17] ), .C(\L2[17] ), .D(\L3[17] ), 
        .Y(Y[17]) );
  NAND3_56 Nand3_1_18 ( .A(S0), .B(n24), .C(inv_R2[18]), .Y(\L0[18] ) );
  NAND3_55 Nand3_2_18 ( .A(n46), .B(n24), .C(R2[18]), .Y(\L1[18] ) );
  NAND3_54 Nand3_3_18 ( .A(n43), .B(R1[18]), .C(inv_R2[18]), .Y(\L2[18] ) );
  NAND3_53 Nand3_4_18 ( .A(n40), .B(R1[18]), .C(R2[18]), .Y(\L3[18] ) );
  NAND4_14 Nand4_0_18 ( .A(\L0[18] ), .B(\L1[18] ), .C(\L2[18] ), .D(\L3[18] ), 
        .Y(Y[18]) );
  NAND3_52 Nand3_1_19 ( .A(S0), .B(n25), .C(inv_R2[19]), .Y(\L0[19] ) );
  NAND3_51 Nand3_2_19 ( .A(n46), .B(n25), .C(R2[19]), .Y(\L1[19] ) );
  NAND3_50 Nand3_3_19 ( .A(n43), .B(R1[19]), .C(inv_R2[19]), .Y(\L2[19] ) );
  NAND3_49 Nand3_4_19 ( .A(n40), .B(R1[19]), .C(R2[19]), .Y(\L3[19] ) );
  NAND4_13 Nand4_0_19 ( .A(\L0[19] ), .B(\L1[19] ), .C(\L2[19] ), .D(\L3[19] ), 
        .Y(Y[19]) );
  NAND3_48 Nand3_1_20 ( .A(S0), .B(n26), .C(inv_R2[20]), .Y(\L0[20] ) );
  NAND3_47 Nand3_2_20 ( .A(n46), .B(n26), .C(R2[20]), .Y(\L1[20] ) );
  NAND3_46 Nand3_3_20 ( .A(n43), .B(R1[20]), .C(inv_R2[20]), .Y(\L2[20] ) );
  NAND3_45 Nand3_4_20 ( .A(n40), .B(R1[20]), .C(R2[20]), .Y(\L3[20] ) );
  NAND4_12 Nand4_0_20 ( .A(\L0[20] ), .B(\L1[20] ), .C(\L2[20] ), .D(\L3[20] ), 
        .Y(Y[20]) );
  NAND3_44 Nand3_1_21 ( .A(S0), .B(n27), .C(inv_R2[21]), .Y(\L0[21] ) );
  NAND3_43 Nand3_2_21 ( .A(n46), .B(n27), .C(R2[21]), .Y(\L1[21] ) );
  NAND3_42 Nand3_3_21 ( .A(n43), .B(R1[21]), .C(inv_R2[21]), .Y(\L2[21] ) );
  NAND3_41 Nand3_4_21 ( .A(n40), .B(R1[21]), .C(R2[21]), .Y(\L3[21] ) );
  NAND4_11 Nand4_0_21 ( .A(\L0[21] ), .B(\L1[21] ), .C(\L2[21] ), .D(\L3[21] ), 
        .Y(Y[21]) );
  NAND3_40 Nand3_1_22 ( .A(S0), .B(n28), .C(inv_R2[22]), .Y(\L0[22] ) );
  NAND3_39 Nand3_2_22 ( .A(n46), .B(n28), .C(R2[22]), .Y(\L1[22] ) );
  NAND3_38 Nand3_3_22 ( .A(n43), .B(R1[22]), .C(inv_R2[22]), .Y(\L2[22] ) );
  NAND3_37 Nand3_4_22 ( .A(n40), .B(R1[22]), .C(R2[22]), .Y(\L3[22] ) );
  NAND4_10 Nand4_0_22 ( .A(\L0[22] ), .B(\L1[22] ), .C(\L2[22] ), .D(\L3[22] ), 
        .Y(Y[22]) );
  NAND3_36 Nand3_1_23 ( .A(S0), .B(n29), .C(inv_R2[23]), .Y(\L0[23] ) );
  NAND3_35 Nand3_2_23 ( .A(n46), .B(n29), .C(R2[23]), .Y(\L1[23] ) );
  NAND3_34 Nand3_3_23 ( .A(n43), .B(R1[23]), .C(inv_R2[23]), .Y(\L2[23] ) );
  NAND3_33 Nand3_4_23 ( .A(n40), .B(R1[23]), .C(R2[23]), .Y(\L3[23] ) );
  NAND4_9 Nand4_0_23 ( .A(\L0[23] ), .B(\L1[23] ), .C(\L2[23] ), .D(\L3[23] ), 
        .Y(Y[23]) );
  NAND3_32 Nand3_1_24 ( .A(S0), .B(n30), .C(inv_R2[24]), .Y(\L0[24] ) );
  NAND3_31 Nand3_2_24 ( .A(n46), .B(n30), .C(R2[24]), .Y(\L1[24] ) );
  NAND3_30 Nand3_3_24 ( .A(n43), .B(R1[24]), .C(inv_R2[24]), .Y(\L2[24] ) );
  NAND3_29 Nand3_4_24 ( .A(n40), .B(R1[24]), .C(R2[24]), .Y(\L3[24] ) );
  NAND4_8 Nand4_0_24 ( .A(\L0[24] ), .B(\L1[24] ), .C(\L2[24] ), .D(\L3[24] ), 
        .Y(Y[24]) );
  NAND3_28 Nand3_1_25 ( .A(S0), .B(n31), .C(inv_R2[25]), .Y(\L0[25] ) );
  NAND3_27 Nand3_2_25 ( .A(n46), .B(n31), .C(R2[25]), .Y(\L1[25] ) );
  NAND3_26 Nand3_3_25 ( .A(n43), .B(R1[25]), .C(inv_R2[25]), .Y(\L2[25] ) );
  NAND3_25 Nand3_4_25 ( .A(n40), .B(R1[25]), .C(R2[25]), .Y(\L3[25] ) );
  NAND4_7 Nand4_0_25 ( .A(\L0[25] ), .B(\L1[25] ), .C(\L2[25] ), .D(\L3[25] ), 
        .Y(Y[25]) );
  NAND3_24 Nand3_1_26 ( .A(S0), .B(n32), .C(inv_R2[26]), .Y(\L0[26] ) );
  NAND3_23 Nand3_2_26 ( .A(n46), .B(n32), .C(R2[26]), .Y(\L1[26] ) );
  NAND3_22 Nand3_3_26 ( .A(n43), .B(R1[26]), .C(inv_R2[26]), .Y(\L2[26] ) );
  NAND3_21 Nand3_4_26 ( .A(n40), .B(R1[26]), .C(R2[26]), .Y(\L3[26] ) );
  NAND4_6 Nand4_0_26 ( .A(\L0[26] ), .B(\L1[26] ), .C(\L2[26] ), .D(\L3[26] ), 
        .Y(Y[26]) );
  NAND3_20 Nand3_1_27 ( .A(S0), .B(n33), .C(inv_R2[27]), .Y(\L0[27] ) );
  NAND3_19 Nand3_2_27 ( .A(n46), .B(n33), .C(R2[27]), .Y(\L1[27] ) );
  NAND3_18 Nand3_3_27 ( .A(n43), .B(R1[27]), .C(inv_R2[27]), .Y(\L2[27] ) );
  NAND3_17 Nand3_4_27 ( .A(n40), .B(R1[27]), .C(R2[27]), .Y(\L3[27] ) );
  NAND4_5 Nand4_0_27 ( .A(\L0[27] ), .B(\L1[27] ), .C(\L2[27] ), .D(\L3[27] ), 
        .Y(Y[27]) );
  NAND3_16 Nand3_1_28 ( .A(S0), .B(n34), .C(inv_R2[28]), .Y(\L0[28] ) );
  NAND3_15 Nand3_2_28 ( .A(n46), .B(n34), .C(R2[28]), .Y(\L1[28] ) );
  NAND3_14 Nand3_3_28 ( .A(n43), .B(R1[28]), .C(inv_R2[28]), .Y(\L2[28] ) );
  NAND3_13 Nand3_4_28 ( .A(n40), .B(R1[28]), .C(R2[28]), .Y(\L3[28] ) );
  NAND4_4 Nand4_0_28 ( .A(\L0[28] ), .B(\L1[28] ), .C(\L2[28] ), .D(\L3[28] ), 
        .Y(Y[28]) );
  NAND3_12 Nand3_1_29 ( .A(S0), .B(n35), .C(inv_R2[29]), .Y(\L0[29] ) );
  NAND3_11 Nand3_2_29 ( .A(n46), .B(n35), .C(R2[29]), .Y(\L1[29] ) );
  NAND3_10 Nand3_3_29 ( .A(n43), .B(R1[29]), .C(inv_R2[29]), .Y(\L2[29] ) );
  NAND3_9 Nand3_4_29 ( .A(n40), .B(R1[29]), .C(R2[29]), .Y(\L3[29] ) );
  NAND4_3 Nand4_0_29 ( .A(\L0[29] ), .B(\L1[29] ), .C(\L2[29] ), .D(\L3[29] ), 
        .Y(Y[29]) );
  NAND3_8 Nand3_1_30 ( .A(S0), .B(n36), .C(inv_R2[30]), .Y(\L0[30] ) );
  NAND3_7 Nand3_2_30 ( .A(n46), .B(n36), .C(R2[30]), .Y(\L1[30] ) );
  NAND3_6 Nand3_3_30 ( .A(n43), .B(R1[30]), .C(inv_R2[30]), .Y(\L2[30] ) );
  NAND3_5 Nand3_4_30 ( .A(n40), .B(R1[30]), .C(R2[30]), .Y(\L3[30] ) );
  NAND4_2 Nand4_0_30 ( .A(\L0[30] ), .B(\L1[30] ), .C(\L2[30] ), .D(\L3[30] ), 
        .Y(Y[30]) );
  NAND3_4 Nand3_1_31 ( .A(S0), .B(n37), .C(inv_R2[31]), .Y(\L0[31] ) );
  NAND3_3 Nand3_2_31 ( .A(n46), .B(n37), .C(R2[31]), .Y(\L1[31] ) );
  NAND3_2 Nand3_3_31 ( .A(n43), .B(R1[31]), .C(inv_R2[31]), .Y(\L2[31] ) );
  NAND3_1 Nand3_4_31 ( .A(n40), .B(R1[31]), .C(R2[31]), .Y(\L3[31] ) );
  NAND4_1 Nand4_0_31 ( .A(\L0[31] ), .B(\L1[31] ), .C(\L2[31] ), .D(\L3[31] ), 
        .Y(Y[31]) );
  INV_X1 U1 ( .A(R2[31]), .ZN(inv_R2[31]) );
  INV_X1 U2 ( .A(R1[31]), .ZN(n37) );
  INV_X1 U3 ( .A(R2[30]), .ZN(inv_R2[30]) );
  INV_X1 U4 ( .A(R1[30]), .ZN(n36) );
  INV_X1 U5 ( .A(R2[29]), .ZN(inv_R2[29]) );
  INV_X1 U6 ( .A(R1[29]), .ZN(n35) );
  INV_X1 U7 ( .A(R2[28]), .ZN(inv_R2[28]) );
  INV_X1 U8 ( .A(R1[28]), .ZN(n34) );
  INV_X1 U9 ( .A(R2[27]), .ZN(inv_R2[27]) );
  INV_X1 U10 ( .A(R1[27]), .ZN(n33) );
  INV_X1 U11 ( .A(R2[26]), .ZN(inv_R2[26]) );
  INV_X1 U12 ( .A(R1[26]), .ZN(n32) );
  INV_X1 U13 ( .A(R2[25]), .ZN(inv_R2[25]) );
  INV_X1 U14 ( .A(R1[25]), .ZN(n31) );
  INV_X1 U15 ( .A(R2[24]), .ZN(inv_R2[24]) );
  INV_X1 U16 ( .A(R1[24]), .ZN(n30) );
  INV_X1 U17 ( .A(R2[23]), .ZN(inv_R2[23]) );
  INV_X1 U18 ( .A(R1[23]), .ZN(n29) );
  INV_X1 U19 ( .A(R2[22]), .ZN(inv_R2[22]) );
  INV_X1 U20 ( .A(R1[22]), .ZN(n28) );
  INV_X1 U21 ( .A(R2[21]), .ZN(inv_R2[21]) );
  INV_X1 U22 ( .A(R1[21]), .ZN(n27) );
  INV_X1 U23 ( .A(R2[20]), .ZN(inv_R2[20]) );
  INV_X1 U24 ( .A(R1[20]), .ZN(n26) );
  INV_X1 U25 ( .A(R2[19]), .ZN(inv_R2[19]) );
  INV_X1 U26 ( .A(R1[19]), .ZN(n25) );
  INV_X1 U27 ( .A(R2[18]), .ZN(inv_R2[18]) );
  INV_X1 U28 ( .A(R1[18]), .ZN(n24) );
  INV_X1 U29 ( .A(R2[17]), .ZN(inv_R2[17]) );
  INV_X1 U30 ( .A(R1[17]), .ZN(n23) );
  INV_X1 U31 ( .A(R2[16]), .ZN(inv_R2[16]) );
  INV_X1 U32 ( .A(R1[16]), .ZN(n22) );
  INV_X1 U33 ( .A(R2[15]), .ZN(inv_R2[15]) );
  INV_X1 U34 ( .A(R2[14]), .ZN(inv_R2[14]) );
  INV_X1 U35 ( .A(R2[13]), .ZN(inv_R2[13]) );
  INV_X1 U36 ( .A(R2[12]), .ZN(inv_R2[12]) );
  INV_X1 U37 ( .A(R2[11]), .ZN(inv_R2[11]) );
  INV_X1 U38 ( .A(R2[10]), .ZN(inv_R2[10]) );
  INV_X1 U39 ( .A(R2[9]), .ZN(inv_R2[9]) );
  INV_X1 U40 ( .A(R2[8]), .ZN(inv_R2[8]) );
  INV_X1 U41 ( .A(R2[7]), .ZN(inv_R2[7]) );
  INV_X1 U42 ( .A(R2[6]), .ZN(inv_R2[6]) );
  INV_X1 U43 ( .A(R2[5]), .ZN(inv_R2[5]) );
  INV_X1 U44 ( .A(R2[0]), .ZN(n194) );
  INV_X1 U45 ( .A(R2[1]), .ZN(n195) );
  INV_X1 U46 ( .A(R2[2]), .ZN(n196) );
  INV_X1 U47 ( .A(R2[3]), .ZN(n197) );
  INV_X1 U48 ( .A(R2[4]), .ZN(n198) );
  INV_X1 U49 ( .A(R1[0]), .ZN(n199) );
  INV_X1 U50 ( .A(R1[1]), .ZN(n200) );
  INV_X1 U51 ( .A(R1[2]), .ZN(n201) );
  INV_X1 U52 ( .A(R1[3]), .ZN(n202) );
  INV_X1 U53 ( .A(R1[4]), .ZN(n203) );
  INV_X1 U54 ( .A(R1[5]), .ZN(n204) );
  INV_X1 U55 ( .A(R1[6]), .ZN(n205) );
  INV_X1 U56 ( .A(R1[7]), .ZN(n206) );
  INV_X1 U57 ( .A(R1[8]), .ZN(n207) );
  INV_X1 U58 ( .A(R1[9]), .ZN(n208) );
  INV_X1 U59 ( .A(R1[10]), .ZN(n209) );
  INV_X1 U60 ( .A(R1[11]), .ZN(n210) );
  INV_X1 U61 ( .A(R1[12]), .ZN(n211) );
  INV_X1 U62 ( .A(R1[13]), .ZN(n212) );
  INV_X1 U63 ( .A(R1[14]), .ZN(n213) );
  INV_X1 U64 ( .A(R1[15]), .ZN(n214) );
endmodule


module DRAM_MEM_DEPTH80_D_SIZE32 ( RESET, CLK, DATAIN, ENABLE, WR_enable, Addr, 
        Dout );
  input [31:0] DATAIN;
  input [31:0] Addr;
  output [31:0] Dout;
  input RESET, CLK, ENABLE, WR_enable;
  wire   n4083, n4085, n4087, n4089, n4091, n4093, n4095, n4097, n4099, n4101,
         n4103, n4105, n4107, n4109, n4111, n4113, n4115, n4117, n4119, n4121,
         n4123, n4125, n4127, n4129, n4131, n4133, n4135, n4137, n4139, n4141,
         n4143, n4145, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n6368, n6369, n6370, n6372, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6407, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6442, n6445, n6448, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6483, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, net253551, net253552, net253553, net253554, net253555,
         net253556, net253557, net253558, net253559, net253560, net253561,
         net253562, net253563, net253564, net253565, net253566, net253567,
         net253568, net253569, net253570, net253571, net253572, net253573,
         net253574, net253575, net253576, net253577, net253578, net253579,
         net253580, net253581, net253582, net253583, net253584, net253585,
         net253586, net253587, net253588, net253589, net253590, net253591,
         net253592, net253593, net253594, net253595, net253596, net253597,
         net253598, net253599, net253600, net253601, net253602, net253603,
         net253604, net253605, net253606, net253607, net253608, net253609,
         net253610, net253611, net253612, net253613, net253614, net253615,
         net253616, net253617, net253618, net253619, net253620, net253621,
         net253622, net253623, net253624, net253625, net253626, net253627,
         net253628, net253629, net253630, net253631, net253632, net253633,
         net253634, net253635, net253636, net253637, net253638, net253639,
         net253640, net253641, net253642, net253643, net253644, net253645,
         net253646, net253647, net253648, net253649, net253650, net253651,
         net253652, net253653, net253654, net253655, net253656, net253657,
         net253658, net253659, net253660, net253661, net253662, net253663,
         net253664, net253665, net253666, net253667, net253668, net253669,
         net253670, net253671, net253672, net253673, net253674, net253675,
         net253676, net253677, net253678, net253679, net253680, net253681,
         net253682, net253683, net253684, net253685, net253686, net253687,
         net253688, net253689, net253690, net253691, net253692, net253693,
         net253694, net253695, net253696, net253697, net253698, net253699,
         net253700, net253701, net253702, net253703, net253704, net253705,
         net253706, net253707, net253708, net253709, net253710, net253711,
         net253712, net253713, net253714, net253715, net253716, net253717,
         net253718, net253719, net253720, net253721, net253722, net253723,
         net253724, net253725, net253726, net253727, net253728, net253729,
         net253730, net253731, net253732, net253733, net253734, net253735,
         net253736, net253737, net253738, net253739, net253740, net253741,
         net253742, net253743, net253744, net253745, net253746, net253747,
         net253748, net253749, net253750, net253751, net253752, net253753,
         net253754, net253755, net253756, net253757, net253758, net253759,
         net253760, net253761, net253762, net253763, net253764, net253765,
         net253766, net253767, net253768, net253769, net253770, net253771,
         net253772, net253773, net253774, net253775, net253776, net253777,
         net253778, net253779, net253780, net253781, net253782, net253783,
         net253784, net253785, net253786, net253787, net253788, net253789,
         net253790, net253791, net253792, net253793, net253794, net253795,
         net253796, net253797, net253798, net253799, net253800, net253801,
         net253802, net253803, net253804, net253805, net253806, net253807,
         net253808, net253809, net253810, net253811, net253812, net253813,
         net253814, net253815, net253816, net253817, net253818, net253819,
         net253820, net253821, net253822, net253823, net253824, net253825,
         net253826, net253827, net253828, net253829, net253830, net253831,
         net253832, net253833, net253834, net253835, net253836, net253837,
         net253838, net253839, net253840, net253841, net253842, net253843,
         net253844, net253845, net253846, net253847, net253848, net253849,
         net253850, net253851, net253852, net253853, net253854, net253855,
         net253856, net253857, net253858, net253859, net253860, net253861,
         net253862, net253863, net253864, net253865, net253866, net253867,
         net253868, net253869, net253870, net253871, net253872, net253873,
         net253874, net253875, net253876, net253877, net253878, net253879,
         net253880, net253881, net253882, net253883, net253884, net253885,
         net253886, net253887, net253888, net253889, net253890, net253891,
         net253892, net253893, net253894, net253895, net253896, net253897,
         net253898, net253899, net253900, net253901, net253902, net253903,
         net253904, net253905, net253906, net253907, net253908, net253909,
         net253910, net253911, net253912, net253913, net253914, net253915,
         net253916, net253917, net253918, net253919, net253920, net253921,
         net253922, net253923, net253924, net253925, net253926, net253927,
         net253928, net253929, net253930, net253931, net253932, net253933,
         net253934, net253935, net253936, net253937, net253938, net253939,
         net253940, net253941, net253942, net253943, net253944, net253945,
         net253946, net253947, net253948, net253949, net253950, net253951,
         net253952, net253953, net253954, net253955, net253956, net253957,
         net253958, net253959, net253960, net253961, net253962, net253963,
         net253964, net253965, net253966, net253967, net253968, net253969,
         net253970, net253971, net253972, net253973, net253974, net253975,
         net253976, net253977, net253978, net253979, net253980, net253981,
         net253982, net253983, net253984, net253985, net253986, net253987,
         net253988, net253989, net253990, net253991, net253992, net253993,
         net253994, net253995, net253996, net253997, net253998, net253999,
         net254000, net254001, net254002, net254003, net254004, net254005,
         net254006, net254007, net254008, net254009, net254010, net254011,
         net254012, net254013, net254014, net254015, net254016, net254017,
         net254018, net254019, net254020, net254021, net254022, net254023,
         net254024, net254025, net254026, net254027, net254028, net254029,
         net254030, net254031, net254032, net254033, net254034, net254035,
         net254036, net254037, net254038, net254039, net254040, net254041,
         net254042, net254043, net254044, net254045, net254046, net254047,
         net254048, net254049, net254050, net254051, net254052, net254053,
         net254054, net254055, net254056, net254057, net254058, net254059,
         net254060, net254061, net254062, net254063, net254064, net254065,
         net254066, net254067, net254068, net254069, net254070, net254071,
         net254072, net254073, net254074, net254075, net254076, net254077,
         net254078, net254079, net254080, net254081, net254082, net254083,
         net254084, net254085, net254086, net254087, net254088, net254089,
         net254090, net254091, net254092, net254093, net254094, net254095,
         net254096, net254097, net254098, net254099, net254100, net254101,
         net254102, net254103, net254104, net254105, net254106, net254107,
         net254108, net254109, net254110, net254111, net254112, net254113,
         net254114, net254115, net254116, net254117, net254118, net254119,
         net254120, net254121, net254122, net254123, net254124, net254125,
         net254126, net254127, net254128, net254129, net254130, net254131,
         net254132, net254133, net254134, net254135, net254136, net254137,
         net254138, net254139, net254140, net254141, net254142, net254143,
         net254144, net254145, net254146, net254147, net254148, net254149,
         net254150, net254151, net254152, net254153, net254154, net254155,
         net254156, net254157, net254158, net254159, net254160, net254161,
         net254162, net254163, net254164, net254165, net254166, net254167,
         net254168, net254169, net254170, net254171, net254172, net254173,
         net254174, net254175, net254176, net254177, net254178, net254179,
         net254180, net254181, net254182, net254183, net254184, net254185,
         net254186, net254187, net254188, net254189, net254190, net254191,
         net254192, net254193, net254194, net254195, net254196, net254197,
         net254198, net254199, net254200, net254201, net254202, net254203,
         net254204, net254205, net254206, net254207, net254208, net254209,
         net254210, net254211, net254212, net254213, net254214, net254215,
         net254216, net254217, net254218, net254219, net254220, net254221,
         net254222, net254223, net254224, net254225, net254226, net254227,
         net254228, net254229, net254230, net254231, net254232, net254233,
         net254234, net254235, net254236, net254237, net254238, net254239,
         net254240, net254241, net254242, net254243, net254244, net254245,
         net254246, net254247, net254248, net254249, net254250, net254251,
         net254252, net254253, net254254, net254255, net254256, net254257,
         net254258, net254259, net254260, net254261, net254262, net254263,
         net254264, net254265, net254266, net254267, net254268, net254269,
         net254270, net254271, net254272, net254273, net254274, net254275,
         net254276, net254277, net254278, net254279, net254280, net254281,
         net254282, net254283, net254284, net254285, net254286, net254287,
         net254288, net254289, net254290, net254291, net254292, net254293,
         net254294, net254295, net254296, net254297, net254298, net254299,
         net254300, net254301, net254302, net254303, net254304, net254305,
         net254306, net254307, net254308, net254309, net254310, net254311,
         net254312, net254313, net254314, net254315, net254316, net254317,
         net254318, n5553, n5555, n5558, n5560, n5604, n5606, n5608, n5610,
         n5646, n5648, n5650, n5652, n5688, n5690, n5692, n5694, n5730, n5732,
         n5734, n5736, n5772, n5774, n5776, n5778, n5814, n5816, n5818, n5820,
         n5856, n5858, n5860, n5862, n5898, n5900, n5902, n5904, n5940, n5942,
         n5944, n5946, n5982, n5984, n5986, n5988, n6024, n6026, n6028, n6030,
         n6066, n6068, n6070, n6072, n6108, n6110, n6112, n6114, n6150, n6152,
         n6154, n6156, n6192, n6194, n6196, n6198, n6234, n6236, n6238, n6240,
         n6276, n6278, n6280, n6282, n6318, n6320, n6322, n6324, n6360, n6362,
         n6364, n6366, n6530, n6532, n6534, n6536, n6572, n6574, n6576, n6578,
         n6614, n6616, n6618, n6620, n6656, n6658, n6660, n6662, n9290, n9292,
         n9294, n9296, n9332, n9334, n9336, n9338, n9374, n9376, n9378, n9380,
         n9416, n9418, n9420, n9422, n9458, n9460, n9462, n9464, n9500, n9502,
         n9504, n9506, n9542, n9544, n9546, n9548, n9602, n9605, n9609, n9613,
         n2676, n2677, n2679, n2681, n2683, n2685, n2687, n2689, n2691, n2693,
         n2695, n2697, n2699, n2701, n2703, n2705, n2707, n2709, n2711, n2713,
         n2715, n2717, n2719, n2721, n2723, n2725, n2727, n2729, n2731, n2733,
         n2735, n2737, n2739, n2740, n2741, n2744, n2776, n2778, n2811, n2812,
         n2815, n2848, n2850, n2883, n2886, n2918, n2921, n2953, n2955, n2988,
         n2990, n3023, n3025, n3058, n3061, n3093, n3096, n3128, n3130, n3163,
         n3165, n3198, n3200, n3233, n3236, n3268, n3270, n3303, n3304, n3306,
         n3339, n3341, n3374, n3376, n3409, n3411, n3444, n3446, n3479, n3481,
         n3514, n3516, n3549, n3551, n3584, n3586, n3619, n3621, n3654, n3656,
         n3689, n3691, n3724, n3726, n3759, n3761, n3794, n3796, n3829, n3831,
         n3864, n3866, n3899, n3901, n3934, n3936, n3969, n3971, n4004, n4006,
         n4039, n4041, n4074, n4076, n4136, n4140, n4176, n4178, n4211, n4213,
         n4246, n4248, n4281, n4283, n4316, n4318, n4351, n4353, n4386, n4388,
         n4421, n4423, n4456, n4458, n4491, n4493, n4526, n4528, n4561, n4563,
         n4596, n4598, n4631, n4633, n4666, n4668, n4701, n4703, n4736, n4738,
         n4771, n4773, n4806, n4808, n4841, n4843, n4876, n4878, n4911, n4913,
         n4946, n4948, n4981, n4983, n5016, n5017, n5019, n5052, n5054, n5087,
         n5089, n5122, n5124, n5157, n5159, n5192, n5194, n5227, n5229, n5262,
         n5264, n5297, n5299, n5332, n5334, n5367, n5369, n5402, n5404, n5437,
         n5439, n5472, n5474, n5507, n5508, n5512, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5554, n5556, n5557, n5559, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5605, n5607, n5609, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5647, n5649,
         n5651, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5689, n5691, n5693, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5731, n5733, n5735, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5773,
         n5775, n5777, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5815, n5817, n5819, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5857, n5859, n5861, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5899, n5901, n5903, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5941, n5943, n5945,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5983, n5985, n5987, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6025, n6027, n6029, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6067, n6069,
         n6071, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6109, n6111, n6113, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6151, n6153, n6155, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6193,
         n6195, n6197, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6235, n6237, n6239, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6277, n6279, n6281, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6319, n6321, n6323, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6361, n6363, n6365,
         n6367, n6371, n6373, n6406, n6408, n6441, n6443, n6444, n6446, n6447,
         n6482, n6484, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6531, n6533, n6535, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6573, n6575, n6577, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6615, n6617,
         n6619, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6657, n6659, n6661, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6674, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9291, n9293, n9295, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9333,
         n9335, n9337, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9375, n9377, n9379, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9417, n9419, n9421, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9459, n9461, n9463, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9501, n9503, n9505,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9543, n9545, n9547, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9603,
         n9604, n9606, n9607, n9608, n9610, n9611, n9612, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n35149, n35150, n35151, n35152,
         n35153, n35154, n35155, n35156, n35157, n35158, n35159, n35160,
         n35161, n35162, n35163, n35164, n35165, n35166, n35167, n35168,
         n35169, n35170, n35171, n35172, n35173, n35174, n35175, n35176,
         n35177, n35178, n35179, n35180, n35181, n35182, n35183, n35184,
         n35185, n35186, n35187, n35188, n35189, n35190, n35191, n35192,
         n35193, n35194, n35195, n35196, n35197, n35198, n35199, n35200,
         n35201, n35202, n35203, n35204, n35205, n35206, n35207, n35208,
         n35209, n35210, n35211, n35212, n35213, n35214, n35215, n35216,
         n35217, n35218, n35219, n35220, n35221, n35222, n35223, n35224,
         n35225, n35226, n35227, n35228, n35229, n35230, n35231, n35232,
         n35233, n35234, n35235, n35236, n35237, n35238, n35239, n35240,
         n35241, n35242, n35243, n35244, n35245, n35246, n35247, n35248,
         n35249, n35250, n35251, n35252, n35253, n35254, n35255, n35256,
         n35257, n35258, n35259, n35260, n35261, n35262, n35263, n35264,
         n35265, n35266, n35267, n35268, n35269, n35270, n35271, n35272,
         n35273, n35274, n35275, n35276, n35277, n35278, n35279, n35280,
         n35281, n35282, n35283, n35284, n35285, n35286, n35287, n35288,
         n35289, n35290, n35291, n35292, n35293, n35294, n35295, n35296,
         n35297, n35298, n35299, n35300, n35301, n35302, n35303, n35304,
         n35305, n35306, n35307, n35308, n35309, n35310, n35311, n35312,
         n35313, n35314, n35315, n35316, n35317, n35318, n35319, n35320,
         n35321, n35322, n35323, n35324, n35325, n35326, n35327, n35328,
         n35329, n35330, n35331, n35332, n35333, n35334, n35335, n35336,
         n35337, n35338, n35339, n35340, n35341, n35342, n35343, n35344,
         n35345, n35346, n35347, n35348, n35349, n35350, n35351, n35352,
         n35353, n35354, n35355, n35356, n35357, n35358, n35359, n35360,
         n35361, n35362, n35363, n35364, n35365, n35366, n35367, n35368,
         n35369, n35370, n35371, n35372, n35373, n35374, n35375, n35376,
         n35377, n35378, n35379, n35380, n35381, n35382, n35383, n35384,
         n35385, n35386, n35387, n35388, n35389, n35390, n35391, n35392,
         n35393, n35394, n35395, n35396, n35397, n35398, n35399, n35400,
         n35401, n35402, n35403, n35404, n35405, n35406, n35407, n35408,
         n35409, n35410, n35411, n35412, n35413, n35414, n35415, n35416,
         n35417, n35418, n35419, n35420, n35421, n35422, n35423, n35424,
         n35425, n35426, n35427, n35428, n35429, n35430, n35431, n35432,
         n35433, n35434, n35435, n35436, n35437, n35438, n35439, n35440,
         n35441, n35442, n35443, n35444, n35445, n35446, n35447, n35448,
         n35449, n35450, n35451, n35452, n35453, n35454, n35455, n35456,
         n35457, n35458, n35459, n35460, n35461, n35462, n35463, n35464,
         n35465, n35466, n35467, n35468, n35469, n35470, n35471, n35472,
         n35473, n35474, n35475, n35476, n35477, n35478, n35479, n35480,
         n35481, n35482, n35483, n35484, n35485, n35486, n35487, n35488,
         n35489, n35490, n35491, n35492, n35493, n35494, n35495, n35496,
         n35497, n35498, n35499, n35500, n35501, n35502, n35503, n35504,
         n35505, n35506, n35507, n35508, n35509, n35510, n35511, n35512,
         n35513, n35514, n35515, n35516, n35517, n35518, n35519, n35520,
         n35521, n35522, n35523, n35524, n35525, n35526, n35527, n35528,
         n35529, n35530, n35531, n35532, n35533, n35534, n35535, n35536,
         n35537, n35538, n35539, n35540, n35541, n35542, n35543, n35544,
         n35545, n35546, n35547, n35548, n35549, n35550, n35551, n35552,
         n35553, n35554, n35555, n35556, n35557, n35558, n35559, n35560,
         n35561, n35562, n35563, n35564, n35565, n35566, n35567, n35568,
         n35569, n35570, n35571, n35572, n35573, n35574, n35575, n35576,
         n35577, n35578, n35579, n35580, n35581, n35582, n35583, n35584,
         n35585, n35586, n35587, n35588, n35589, n35590, n35591, n35592,
         n35593, n35594, n35595, n35596, n35597, n35598, n35599, n35600,
         n35601, n35602, n35603, n35604, n35605, n35606, n35607, n35608,
         n35609, n35610, n35611, n35612, n35613, n35614, n35615, n35616,
         n35617, n35618, n35619, n35620, n35621, n35622, n35623, n35624,
         n35625, n35626, n35627, n35628, n35629, n35630, n35631, n35632,
         n35633, n35634, n35635, n35636, n35637, n35638, n35639, n35640,
         n35641, n35642, n35643, n35644, n35645, n35646, n35647, n35648,
         n35649, n35650, n35651, n35652, n35653, n35654, n35655, n35656,
         n35657, n35658, n35659, n35660, n35661, n35662, n35663, n35664,
         n35665, n35666, n35667, n35668, n35669, n35670, n35671, n35672,
         n35673, n35674, n35675, n35676, n35677, n35678, n35679, n35680,
         n35681, n35682, n35683, n35684, n35685, n35686, n35687, n35688,
         n35689, n35690, n35691, n35692, n35693, n35694, n35695, n35696,
         n35697, n35698, n35699, n35700, n35701, n35702, n35703, n35704,
         n35705, n35706, n35707, n35708, n35709, n35710, n35711, n35712,
         n35713, n35714, n35715, n35716, n35717, n35718, n35719, n35720,
         n35721, n35722, n35723, n35724, n35725, n35726, n35727, n35728,
         n35729, n35730, n35731, n35732, n35733, n35734, n35735, n35736,
         n35737, n35738, n35739, n35740, n35741, n35742, n35743, n35744,
         n35745, n35746, n35747, n35748, n35749, n35750, n35751, n35752,
         n35753, n35754, n35755, n35756, n35757, n35758, n35759, n35760,
         n35761, n35762, n35763, n35764, n35765, n35766, n35767, n35768,
         n35769, n35770, n35771, n35772, n35773, n35774, n35775, n35776,
         n35777, n35778, n35779, n35780, n35781, n35782, n35783, n35784,
         n35785, n35786, n35787, n35788, n35789, n35790, n35791, n35792,
         n35793, n35794, n35795, n35796, n35797, n35798, n35799, n35800,
         n35801, n35802, n35803, n35804, n35805, n35806, n35807, n35808,
         n35809, n35810, n35811, n35812, n35813, n35814, n35815, n35816,
         n35817, n35818, n35819, n35820, n35821, n35822, n35823, n35824,
         n35825, n35826, n35827, n35828, n35829, n35830, n35831, n35832,
         n35833, n35834, n35835, n35836, n35837, n35838, n35839, n35840,
         n35841, n35842, n35843, n35844, n35845, n35846, n35847, n35848,
         n35849, n35850, n35851, n35852, n35853, n35854, n35855, n35856,
         n35857, n35858, n35859, n35860, n35861, n35862, n35863, n35864,
         n35865, n35866, n35867, n35868, n35869, n35870, n35871, n35872,
         n35873, n35874, n35875, n35876, n35877, n35878, n35879, n35880,
         n35881, n35882, n35883, n35884, n35885, n35886, n35887, n35888,
         n35889, n35890, n35891, n35892, n35893, n35894, n35895, n35896,
         n35897, n35898, n35899, n35900, n35901, n35902, n35903, n35904,
         n35905, n35906, n35907, n35908, n35909, n35910, n35911, n35912,
         n35913, n35914, n35915, n35916, n35917, n35918, n35919, n35920,
         n35921, n35922, n35923, n35924, n35925, n35926, n35927, n35928,
         n35929, n35930, n35931, n35932, n35933, n35934, n35935, n35936,
         n35937, n35938, n35939, n35940, n35941, n35942, n35943, n35944,
         n35945, n35946, n35947, n35948, n35949, n35950, n35951, n35952,
         n35953, n35954, n35955, n35956, n35957, n35958, n35959, n35960,
         n35961, n35962, n35963, n35964, n35965, n35966, n35967, n35968,
         n35969, n35970, n35971, n35972, n35973, n35974, n35975, n35976,
         n35977, n35978, n35979, n35980, n35981, n35982, n35983, n35984,
         n35985, n35986, n35987, n35988, n35989, n35990, n35991, n35992,
         n35993, n35994, n35995, n35996, n35997, n35998, n35999, n36000,
         n36001, n36002, n36003, n36004, n36005, n36006, n36007, n36008,
         n36009, n36010, n36011, n36012, n36013, n36014, n36015, n36016,
         n36017, n36018, n36019, n36020, n36021, n36022, n36023, n36024,
         n36025, n36026, n36027, n36028, n36029, n36030, n36031, n36032,
         n36033, n36034, n36035, n36036, n36037, n36038, n36039, n36040,
         n36041, n36042, n36043, n36044, n36045, n36046, n36047, n36048,
         n36049, n36050, n36051, n36052, n36053, n36054, n36055, n36056,
         n36057, n36058, n36059, n36060, n36061, n36062, n36063, n36064,
         n36065, n36066, n36067, n36068, n36069, n36070, n36071, n36072,
         n36073, n36074, n36075, n36076, n36077, n36078, n36079, n36080,
         n36081, n36082, n36083, n36084, n36085, n36086, n36087, n36088,
         n36089, n36090, n36091, n36092, n36093, n36094, n36095, n36096,
         n36097, n36098, n36099, n36100, n36101, n36102, n36103, n36104,
         n36105, n36106, n36107, n36108, n36109, n36110, n36111, n36112,
         n36113, n36114, n36115, n36116, n36117, n36118, n36119, n36120,
         n36121, n36122, n36123, n36124, n36125, n36126, n36127, n36128,
         n36129, n36130, n36131, n36132, n36133, n36134, n36135, n36136,
         n36137, n36138, n36139, n36140, n36141, n36142, n36143, n36144,
         n36145, n36146, n36147, n36148, n36149, n36150, n36151, n36152,
         n36153, n36154, n36155, n36156, n36157, n36158, n36159, n36160,
         n36161, n36162, n36163, n36164, n36165, n36166, n36167, n36168,
         n36169, n36170, n36171, n36172, n36173, n36174, n36175, n36176,
         n36177, n36178, n36179, n36180, n36181, n36182, n36183, n36184,
         n36185, n36186, n36187, n36188, n36189, n36190, n36191, n36192,
         n36193, n36194, n36195, n36196, n36197, n36198, n36199, n36200,
         n36201, n36202, n36203, n36204, n36205, n36206, n36207, n36208,
         n36209, n36210, n36211, n36212, n36213, n36214, n36215, n36216,
         n36217, n36218, n36219, n36220, n36221, n36222, n36223, n36224,
         n36225, n36226, n36227, n36228, n36229, n36230, n36231, n36232,
         n36233, n36234, n36235, n36236, n36237, n36238, n36239, n36240,
         n36241, n36242, n36243, n36244, n36245, n36246, n36247, n36248,
         n36249, n36250, n36251, n36252, n36253, n36254, n36255, n36256,
         n36257, n36258, n36259, n36260, n36261, n36262, n36263, n36264,
         n36265, n36266, n36267, n36268, n36269, n36270, n36271, n36272,
         n36273, n36274, n36275, n36276, n36277, n36278, n36279, n36280,
         n36281, n36282, n36283, n36284, n36285, n36286, n36287, n36288,
         n36289, n36290, n36291, n36292, n36293, n36294, n36295, n36296,
         n36297, n36298, n36299, n36300, n36301, n36302, n36303, n36304,
         n36305, n36306, n36307, n36308, n36309, n36310, n36311, n36312,
         n36313, n36314, n36315, n36316, n36317, n36318, n36319, n36320,
         n36321, n36322, n36323, n36324, n36325, n36326, n36327, n36328,
         n36329, n36330, n36331, n36332, n36333, n36334, n36335, n36336,
         n36337, n36338, n36339, n36340, n36341, n36342, n36343, n36344,
         n36345, n36346, n36347, n36348, n36349, n36350, n36351, n36352,
         n36353, n36354, n36355, n36356, n36357, n36358, n36359, n36360,
         n36361, n36362, n36363, n36364, n36365, n36366, n36367, n36368,
         n36369, n36370, n36371, n36372, n36373, n36374, n36375, n36376,
         n36377, n36378, n36379, n36380, n36381, n36382, n36383, n36384,
         n36385, n36386, n36387, n36388, n36389, n36390, n36391, n36392,
         n36393, n36394, n36395, n36396, n36397, n36398, n36399, n36400,
         n36401, n36402, n36403, n36404, n36405, n36406, n36407, n36408,
         n36409, n36410, n36411, n36412, n36413, n36414, n36415, n36416,
         n36417, n36418, n36419, n36420, n36421, n36422, n36423, n36424,
         n36425, n36426, n36427, n36428, n36429, n36430, n36431, n36432,
         n36433, n36434, n36435, n36436, n36437, n36438, n36439, n36440,
         n36441, n36442, n36443, n36444, n36445, n36446, n36447, n36448,
         n36449, n36450, n36451, n36452, n36453, n36454, n36455, n36456,
         n36457, n36458, n36459, n36460, n36461, n36462, n36463, n36464,
         n36465, n36466, n36467, n36468, n36469, n36470, n36471, n36472,
         n36473, n36474, n36475, n36476, n36477, n36478, n36479, n36480,
         n36481, n36482, n36483, n36484, n36485, n36486, n36487, n36488,
         n36489, n36490, n36491, n36492, n36493, n36494, n36495, n36496,
         n36497, n36498, n36499, n36500, n36501, n36502, n36503, n36504,
         n36505, n36506, n36507, n36508, n36509, n36510, n36511, n36512,
         n36513, n36514, n36515, n36516, n36517, n36518, n36519, n36520,
         n36521, n36522, n36523, n36524, n36525, n36526, n36527, n36528,
         n36529, n36530, n36531, n36532, n36533, n36534, n36535, n36536,
         n36537, n36538, n36539, n36540, n36541, n36542, n36543, n36544,
         n36545, n36546, n36547, n36548, n36549, n36550, n36551, n36552,
         n36553, n36554, n36555, n36556, n36557, n36558, n36559, n36560,
         n36561, n36562, n36563, n36564, n36565, n36566, n36567, n36568,
         n36569, n36570, n36571, n36572, n36573, n36574, n36575, n36576,
         n36577, n36578, n36579, n36580, n36581, n36582, n36583, n36584,
         n36585, n36586, n36587, n36588, n36589, n36590, n36591, n36592,
         n36593, n36594, n36595, n36596, n36597, n36598, n36599, n36600,
         n36601, n36602, n36603, n36604, n36605, n36606, n36607, n36608,
         n36609, n36610, n36611, n36612, n36613, n36614, n36615, n36616,
         n36617, n36618, n36619, n36620, n36621, n36622, n36623, n36624,
         n36625, n36626, n36627, n36628, n36629, n36630, n36631, n36632,
         n36633, n36634, n36635, n36636, n36637, n36638, n36639, n36640,
         n36641, n36642, n36643, n36644, n36645, n36646, n36647, n36648,
         n36649, n36650, n36651, n36652, n36653, n36654, n36655, n36656,
         n36657, n36658, n36659, n36660, n36661, n36662, n36663, n36664,
         n36665, n36666, n36667, n36668, n36669, n36670, n36671, n36672,
         n36673, n36674, n36675, n36676, n36677, n36678, n36679, n36680,
         n36681, n36682, n36683, n36684, n36685, n36686, n36687, n36688,
         n36689, n36690, n36691, n36692, n36693, n36694, n36695, n36696,
         n36697, n36698, n36699, n36700, n36701, n36702, n36703, n36704,
         n36705, n36706, n36707, n36708, n36709, n36710, n36711, n36712,
         n36713, n36714, n36715, n36716, n36717, n36718, n36719, n36720,
         n36721, n36722, n36723, n36724, n36725, n36726, n36727, n36728,
         n36729, n36730, n36731, n36732, n36733, n36734, n36735, n36736,
         n36737, n36738, n36739, n36740, n36741, n36742, n36743, n36744,
         n36745, n36746, n36747, n36748, n36749, n36750, n36751, n36752,
         n36753, n36754, n36755, n36756, n36757, n36758, n36759, n36760,
         n36761, n36762, n36763, n36764, n36765, n36766, n36767, n36768,
         n36769, n36770, n36771, n36772, n36773, n36774, n36775, n36776,
         n36777, n36778, n36779, n36780, n36781, n36782, n36783, n36784,
         n36785, n36786, n36787, n36788, n36789, n36790, n36791, n36792,
         n36793, n36794, n36795, n36796, n36797, n36798, n36799, n36800,
         n36801, n36802, n36803, n36804, n36805, n36806, n36807, n36808,
         n36809, n36810, n36811, n36812, n36813, n36814, n36815, n36816,
         n36817, n36818, n36819, n36820, n36821, n36822, n36823, n36824,
         n36825, n36826, n36827, n36828, n36829, n36830, n36831, n36832,
         n36833, n36834, n36835, n36836, n36837, n36838, n36839, n36840,
         n36841, n36842, n36843, n36844, n36845, n36846, n36847, n36848,
         n36849, n36850, n36851, n36852, n36853, n36854, n36855, n36856,
         n36857, n36858, n36859, n36860, n36861, n36862, n36863, n36864,
         n36865, n36866, n36867, n36868, n36869, n36870, n36871, n36872,
         n36873, n36874, n36875, n36876, n36877, n36878, n36879, n36880,
         n36881, n36882, n36883, n36884, n36885, n36886, n36887, n36888,
         n36889, n36890, n36891, n36892, n36893, n36894, n36895, n36896,
         n36897, n36898, n36899, n36900, n36901, n36902, n36903, n36904,
         n36905, n36906, n36907, n36908, n36909, n36910, n36911, n36912,
         n36913, n36914, n36915, n36916, n36917, n36918, n36919, n36920,
         n36921, n36922, n36923, n36924, n36925, n36926, n36927, n36928,
         n36929, n36930, n36931, n36932, n36933, n36934, n36935, n36936,
         n36937, n36938, n36939, n36940, n36941, n36942, n36943, n36944,
         n36945, n36946, n36947, n36948, n36949, n36950, n36951, n36952,
         n36953, n36954, n36955, n36956, n36957, n36958, n36959, n36960,
         n36961, n36962, n36963, n36964, n36965, n36966, n36967, n36968,
         n36969, n36970, n36971, n36972, n36973, n36974, n36975, n36976,
         n36977, n36978, n36979, n36980, n36981, n36982, n36983, n36984,
         n36985, n36986, n36987, n36988, n36989, n36990, n36991, n36992,
         n36993, n36994, n36995, n36996, n36997, n36998, n36999, n37000,
         n37001, n37002, n37003, n37004, n37005, n37006, n37007, n37008,
         n37009, n37010, n37011, n37012, n37013, n37014, n37015, n37016,
         n37017, n37018, n37019, n37020, n37021, n37022, n37023, n37024,
         n37025, n37026, n37027, n37028, n37029, n37030, n37031, n37032,
         n37033, n37034, n37035, n37036, n37037, n37038, n37039, n37040,
         n37041, n37042, n37043, n37044, n37045, n37046, n37047, n37048,
         n37049, n37050, n37051, n37052, n37053, n37054, n37055, n37056,
         n37057, n37058, n37059, n37060, n37061, n37062, n37063, n37064,
         n37065, n37066, n37067, n37068, n37069, n37070, n37071, n37072,
         n37073, n37074, n37075, n37076, n37077, n37078, n37079, n37080,
         n37081, n37082, n37083, n37084, n37085, n37086, n37087, n37088,
         n37089, n37090, n37091, n37092, n37093, n37094, n37095, n37096,
         n37097, n37098, n37099, n37100, n37101, n37102, n37103, n37104,
         n37105, n37106, n37107, n37108, n37109, n37110, n37111, n37112,
         n37113, n37114, n37115, n37116, n37117, n37118, n37119, n37120,
         n37121, n37122, n37123, n37124, n37125, n37126, n37127, n37128,
         n37129, n37130, n37131, n37132, n37133, n37134, n37135, n37136,
         n37137, n37138, n37139, n37140, n37141, n37142, n37143, n37144,
         n37145, n37146, n37147, n37148, n37149, n37150, n37151, n37152,
         n37153, n37154, n37155, n37156, n37157, n37158, n37159, n37160,
         n37161, n37162, n37163, n37164, n37165, n37166, n37167, n37168,
         n37169, n37170, n37171, n37172, n37173, n37174, n37175, n37176,
         n37177, n37178, n37179, n37180, n37181, n37182, n37183, n37184,
         n37185, n37186, n37187, n37188, n37189, n37190, n37191, n37192,
         n37193, n37194, n37195, n37196, n37197, n37198, n37199, n37200,
         n37201, n37202, n37203, n37204, n37205, n37206, n37207, n37208,
         n37209, n37210, n37211, n37212, n37213, n37214, n37215, n37216,
         n37217, n37218, n37219, n37220, n37221, n37222, n37223, n37224,
         n37225, n37226, n37227, n37228, n37229, n37230, n37231, n37232,
         n37233, n37234, n37235, n37236, n37237, n37238, n37239, n37240,
         n37241, n37242, n37243, n37244, n37245, n37246, n37247, n37248,
         n37249, n37250, n37251, n37252, n37253, n37254, n37255, n37256,
         n37257, n37258, n37259, n37260, n37261, n37262, n37263, n37264,
         n37265, n37266, n37267, n37268, n37269, n37270, n37271, n37272,
         n37273, n37274, n37275, n37276, n37277, n37278, n37279, n37280,
         n37281, n37282, n37283, n37284, n37285, n37286, n37287, n37288,
         n37289, n37290, n37291, n37292, n37293, n37294, n37295, n37296,
         n37297, n37298, n37299, n37300, n37301, n37302, n37303, n37304,
         n37305, n37306, n37307, n37308, n37309, n37310, n37311, n37312,
         n37313, n37314, n37315, n37316, n37317, n37318, n37319, n37320,
         n37321, n37322, n37323, n37324, n37325, n37326, n37327, n37328,
         n37329, n37330, n37331, n37332, n37333, n37334, n37335, n37336,
         n37337, n37338, n37339, n37340, n37341, n37342, n37343, n37344,
         n37345, n37346, n37347, n37348, n37349, n37350, n37351, n37352,
         n37353, n37354, n37355, n37356, n37357, n37358, n37359, n37360,
         n37361, n37362, n37363, n37364, n37365, n37366, n37367, n37368,
         n37369, n37370, n37371, n37372, n37373, n37374, n37375, n37376,
         n37377, n37378, n37379, n37380, n37381, n37382, n37383, n37384,
         n37385, n37386, n37387, n37388, n37389, n37390, n37391, n37392,
         n37393, n37394, n37395, n37396, n37397, n37398, n37399, n37400,
         n37401, n37402, n37403, n37404, n37405, n37406, n37407, n37408,
         n37409, n37410, n37411, n37412, n37413, n37414, n37415, n37416,
         n37417, n37418, n37419, n37420, n37421, n37422, n37423, n37424,
         n37425, n37426, n37427, n37428, n37429, n37430, n37431, n37432,
         n37433, n37434, n37435, n37436, n37437, n37438, n37439, n37440,
         n37441, n37442, n37443, n37444, n37445, n37446, n37447, n37448,
         n37449, n37450, n37451, n37452, n37453, n37454, n37455, n37456,
         n37457, n37458, n37459, n37460, n37461, n37462, n37463, n37464,
         n37465, n37466, n37467, n37468, n37469, n37470, n37471, n37472,
         n37473, n37474, n37475, n37476, n37477, n37478, n37479, n37480,
         n37481, n37482, n37483, n37484, n37485, n37486, n37487, n37488,
         n37489, n37490, n37491, n37492, n37493, n37494, n37495, n37496,
         n37497, n37498, n37499, n37500, n37501, n37502, n37503, n37504,
         n37505, n37506, n37507, n37508, n37509, n37510, n37511, n37512,
         n37513, n37514, n37515, n37516, n37517, n37518, n37519, n37520,
         n37521, n37522, n37523, n37524, n37525, n37526, n37527, n37528,
         n37529, n37530, n37531, n37532, n37533, n37534, n37535, n37536,
         n37537, n37538, n37539, n37540, n37541, n37542, n37543, n37544,
         n37545, n37546, n37547, n37548, n37549, n37550, n37551, n37552,
         n37553, n37554, n37555, n37556, n37557, n37558, n37559, n37560,
         n37561, n37562, n37563, n37564, n37565, n37566, n37567, n37568,
         n37569, n37570, n37571, n37572, n37573, n37574, n37575, n37576,
         n37577, n37578, n37579, n37580, n37581, n37582, n37583, n37584,
         n37585, n37586, n37587, n37588, n37589, n37590, n37591, n37592,
         n37593, n37594, n37595, n37596, n37597, n37598, n37599, n37600,
         n37601, n37602, n37603, n37604, n37605, n37606, n37607, n37608,
         n37609, n37610, n37611, n37612, n37613, n37614, n37615, n37616,
         n37617, n37618, n37619, n37620, n37621, n37622, n37623, n37624,
         n37625, n37626, n37627, n37628, n37629, n37630, n37631, n37632,
         n37633, n37634, n37635, n37636, n37637, n37638, n37639, n37640,
         n37641, n37642, n37643, n37644, n37645, n37646, n37647, n37648,
         n37649, n37650, n37651, n37652, n37653, n37654, n37655, n37656,
         n37657, n37658, n37659, n37660, n37661, n37662, n37663, n37664,
         n37665, n37666, n37667, n37668, n37669, n37670, n37671, n37672,
         n37673, n37674, n37675, n37676, n37677, n37678, n37679, n37680,
         n37681, n37682, n37683, n37684, n37685, n37686, n37687, n37688,
         n37689, n37690, n37691, n37692, n37693, n37694, n37695, n37696,
         n37697, n37698, n37699, n37700, n37701, n37702, n37703, n37704,
         n37705, n37706, n37707, n37708, n37709, n37710, n37711, n37712,
         n37713, n37714, n37715, n37716, n37717, n37718, n37719, n37720,
         n37721, n37722, n37723, n37724, n37725, n37726, n37727, n37728,
         n37729, n37730, n37731, n37732, n37733, n37734, n37735, n37736,
         n37737, n37738, n37739, n37740, n37741, n37742, n37743, n37744,
         n37745, n37746, n37747, n37748, n37749, n37750, n37751, n37752,
         n37753, n37754, n37755, n37756, n37757, n37758, n37759, n37760,
         n37761, n37762, n37763, n37764, n37765, n37766, n37767, n37768,
         n37769, n37770, n37771, n37772, n37773, n37774, n37775, n37776,
         n37777, n37778, n37779, n37780, n37781, n37782, n37783, n37784,
         n37785, n37786, n37787, n37788, n37789, n37790, n37791, n37792,
         n37793, n37794, n37795, n37796, n37797, n37798, n37799, n37800,
         n37801, n37802, n37803, n37804, n37805, n37806, n37807, n37808,
         n37809, n37810, n37811, n37812, n37813, n37814, n37815, n37816,
         n37817, n37818, n37819, n37820, n37821, n37822, n37823, n37824,
         n37825, n37826, n37827, n37828, n37829, n37830, n37831, n37832,
         n37833, n37834, n37835, n37836, n37837, n37838, n37839, n37840,
         n37841, n37842, n37843, n37844, n37845, n37846, n37847, n37848,
         n37849, n37850, n37851, n37852, n37853, n37854, n37855, n37856,
         n37857, n37858, n37859, n37860, n37861, n37862, n37863, n37864,
         n37865, n37866, n37867, n37868, n37869, n37870, n37871, n37872,
         n37873, n37874, n37875, n37876, n37877, n37878, n37879, n37880,
         n37881, n37882, n37883, n37884, n37885, n37886, n37887, n37888,
         n37889, n37890, n37891, n37892, n37893, n37894, n37895, n37896,
         n37897, n37898, n37899, n37900, n37901, n37902, n37903, n37904,
         n37905, n37906, n37907, n37908, n37909, n37910, n37911, n37912,
         n37913, n37914, n37915, n37916, n37917, n37918, n37919, n37920,
         n37921, n37922, n37923, n37924, n37925, n37926, n37927, n37928,
         n37929, n37930, n37931, n37932, n37933, n37934, n37935, n37936,
         n37937, n37938, n37939, n37940, n37941, n37942, n37943, n37944,
         n37945, n37946, n37947, n37948, n37949, n37950, n37951, n37952,
         n37953, n37954, n37955, n37956, n37957, n37958, n37959, n37960,
         n37961, n37962, n37963, n37964, n37965, n37966, n37967, n37968,
         n37969, n37970, n37971, n37972, n37973, n37974, n37975, n37976,
         n37977, n37978, n37979, n37980, n37981, n37982, n37983, n37984,
         n37985, n37986, n37987, n37988, n37989, n37990, n37991, n37992,
         n37993, n37994, n37995, n37996, n37997, n37998, n37999, n38000,
         n38001, n38002, n38003, n38004, n38005, n38006, n38007, n38008,
         n38009, n38010, n38011, n38012, n38013, n38014, n38015, n38016,
         n38017, n38018, n38019, n38020, n38021, n38022, n38023, n38024,
         n38025, n38026, n38027, n38028, n38029, n38030, n38031, n38032,
         n38033, n38034, n38035, n38036, n38037, n38038, n38039, n38040,
         n38041, n38042, n38043, n38044, n38045, n38046, n38047, n38048,
         n38049, n38050, n38051, n38052, n38053, n38054, n38055, n38056,
         n38057, n38058, n38059, n38060, n38061, n38062, n38063, n38064,
         n38065, n38066, n38067, n38068, n38069, n38070, n38071, n38072,
         n38073, n38074, n38075, n38076, n38077, n38078, n38079, n38080,
         n38081, n38082, n38083, n38084, n38085, n38086, n38087, n38088,
         n38089, n38090, n38091, n38092, n38093, n38094, n38095, n38096,
         n38097, n38098, n38099, n38100, n38101, n38102, n38103, n38104,
         n38105, n38106, n38107, n38108, n38109, n38110, n38111, n38112,
         n38113, n38114, n38115, n38116, n38117, n38118, n38119, n38120,
         n38121, n38122, n38123, n38124, n38125, n38126, n38127, n38128,
         n38129, n38130, n38131, n38132, n38133, n38134, n38135, n38136,
         n38137, n38138, n38139, n38140, n38141, n38142, n38143, n38144,
         n38145, n38146, n38147, n38148, n38149, n38150, n38151, n38152,
         n38153, n38154, n38155, n38156, n38157, n38158, n38159, n38160,
         n38161, n38162, n38163, n38164, n38165, n38166, n38167, n38168,
         n38169, n38170, n38171, n38172, n38173, n38174, n38175, n38176,
         n38177, n38178, n38179, n38180, n38181, n38182, n38183, n38184,
         n38185, n38186, n38187, n38188, n38189, n38190, n38191, n38192,
         n38193, n38194, n38195, n38196, n38197, n38198, n38199, n38200,
         n38201, n38202, n38203, n38204, n38205, n38206, n38207, n38208,
         n38209, n38210, n38211, n38212, n38213, n38214, n38215, n38216,
         n38217, n38218, n38219, n38220, n38221, n38222, n38223, n38224,
         n38225, n38226, n38227, n38228, n38229, n38230, n38231, n38232,
         n38233, n38234, n38235, n38236, n38237, n38238, n38239, n38240,
         n38241, n38242, n38243, n38244, n38245, n38246, n38247, n38248,
         n38249, n38250, n38251, n38252, n38253, n38254, n38255, n38256,
         n38257, n38258, n38259, n38260, n38261, n38262, n38263, n38264,
         n38265, n38266, n38267, n38268, n38269, n38270, n38271, n38272,
         n38273, n38274, n38275, n38276, n38277, n38278, n38279, n38280,
         n38281, n38282, n38283, n38284, n38285, n38286, n38287, n38288,
         n38289, n38290, n38291, n38292, n38293, n38294, n38295, n38296,
         n38297, n38298, n38299, n38300, n38301, n38302, n38303, n38304,
         n38305, n38306, n38307, n38308, n38309, n38310, n38311, n38312,
         n38313, n38314, n38315, n38316, n38317, n38318, n38319, n38320,
         n38321, n38322, n38323, n38324, n38325, n38326, n38327, n38328,
         n38329, n38330, n38331, n38332, n38333, n38334, n38335, n38336,
         n38337, n38338, n38339, n38340, n38341, n38342, n38343, n38344,
         n38345, n38346, n38347, n38348, n38349, n38350, n38351, n38352,
         n38353, n38354, n38355, n38356, n38357, n38358, n38359, n38360,
         n38361, n38362, n38363, n38364, n38365, n38366, n38367, n38368,
         n38369, n38370, n38371, n38372, n38373, n38374, n38375, n38376,
         n38377, n38378, n38379, n38380, n38381, n38382, n38383, n38384,
         n38385, n38386, n38387, n38388, n38389, n38390, n38391, n38392,
         n38393, n38394, n38395, n38396, n38397, n38398, n38399, n38400,
         n38401, n38402, n38403, n38404, n38405, n38406, n38407, n38408,
         n38409, n38410, n38411, n38412, n38413, n38414, n38415, n38416,
         n38417, n38418, n38419, n38420, n38421, n38422, n38423, n38424,
         n38425, n38426, n38427, n38428, n38429, n38430, n38431, n38432,
         n38433, n38434, n38435, n38436, n38437, n38438, n38439, n38440,
         n38441, n38442, n38443, n38444, n38445, n38446, n38447, n38448,
         n38449, n38450, n38451, n38452, n38453, n38454, n38455, n38456,
         n38457, n38458, n38459, n38460, n38461, n38462, n38463, n38464,
         n38465, n38466, n38467, n38468, n38469, n38470, n38471, n38472,
         n38473, n38474, n38475, n38476, n38477, n38478, n38479, n38480,
         n38481, n38482, n38483, n38484, n38485, n38486, n38487, n38488,
         n38489, n38490, n38491, n38492, n38493, n38494, n38495, n38496,
         n38497, n38498, n38499, n38500, n38501, n38502, n38503, n38504,
         n38505, n38506, n38507, n38508, n38509, n38510, n38511, n38512,
         n38513, n38514, n38515, n38516, n38517, n38518, n38519, n38520,
         n38521, n38522, n38523, n38524, n38525, n38526, n38527, n38528,
         n38529, n38530, n38531, n38532, n38533, n38534, n38535, n38536,
         n38537, n38538, n38539, n38540, n38541, n38542, n38543, n38544,
         n38545, n38546, n38547, n38548, n38549, n38550, n38551, n38552,
         n38553, n38554, n38555, n38556, n38557, n38558, n38559, n38560,
         n38561, n38562, n38563, n38564, n38565, n38566, n38567, n38568,
         n38569, n38570, n38571, n38572, n38573, n38574, n38575, n38576,
         n38577, n38578, n38579, n38580, n38581, n38582, n38583, n38584,
         n38585, n38586, n38587, n38588, n38589, n38590, n38591, n38592,
         n38593, n38594, n38595, n38596, n38597, n38598, n38599, n38600,
         n38601, n38602, n38603, n38604, n38605, n38606, n38607, n38608,
         n38609, n38610, n38611, n38612, n38613, n38614, n38615, n38616,
         n38617, n38618, n38619, n38620, n38621, n38622, n38623, n38624,
         n38625, n38626, n38627, n38628, n38629, n38630, n38631, n38632,
         n38633, n38634, n38635, n38636, n38637, n38638, n38639, n38640,
         n38641, n38642, n38643, n38644, n38645, n38646, n38647, n38648,
         n38649, n38650, n38651, n38652, n38653, n38654, n38655, n38656,
         n38657, n38658, n38659, n38660, n38661, n38662, n38663, n38664,
         n38665, n38666, n38667, n38668, n38669, n38670, n38671, n38672,
         n38673, n38674, n38675, n38676, n38677, n38678, n38679, n38680,
         n38681, n38682, n38683, n38684, n38685, n38686, n38687, n38688,
         n38689, n38690, n38691, n38692, n38693, n38694, n38695, n38696,
         n38697, n38698, n38699, n38700, n38701, n38702, n38703, n38704,
         n38705, n38706, n38707, n38708, n38709, n38710, n38711, n38712,
         n38713, n38714, n38715, n38716, n38717, n38718, n38719, n38720,
         n38721, n38722, n38723, n38724, n38725, n38726, n38727, n38728,
         n38729, n38730, n38731, n38732, n38733, n38734, n38735, n38736,
         n38737, n38738, n38739, n38740, n38741, n38742, n38743, n38744,
         n38745, n38746, n38747, n38748, n38749, n38750, n38751, n38752,
         n38753, n38754, n38755, n38756, n38757, n38758, n38759, n38760,
         n38761, n38762, n38763, n38764, n38765, n38766, n38767, n38768,
         n38769, n38770, n38771, n38772, n38773, n38774, n38775, n38776,
         n38777, n38778, n38779, n38780, n38781, n38782, n38783, n38784,
         n38785, n38786, n38787, n38788, n38789, n38790, n38791, n38792,
         n38793, n38794, n38795, n38796, n38797, n38798, n38799, n38800,
         n38801, n38802, n38803, n38804, n38805, n38806, n38807, n38808,
         n38809, n38810, n38811, n38812, n38813, n38814, n38815, n38816,
         n38817, n38818, n38819, n38820, n38821, n38822, n38823, n38824,
         n38825, n38826, n38827, n38828, n38829, n38830, n38831, n38832,
         n38833, n38834, n38835, n38836, n38837, n38838, n38839, n38840,
         n38841, n38842, n38843, n38844, n38845, n38846, n38847, n38848,
         n38849, n38850, n38851, n38852, n38853, n38854, n38855, n38856,
         n38857, n38858, n38859, n38860, n38861, n38862, n38863, n38864,
         n38865, n38866, n38867, n38868, n38869, n38870, n38871, n38872,
         n38873, n38874, n38875, n38876, n38877, n38878, n38879, n38880,
         n38881, n38882, n38883, n38884, n38885, n38886, n38887, n38888,
         n38889, n38890, n38891, n38892, n38893, n38894, n38895, n38896,
         n38897, n38898, n38899, n38900, n38901, n38902, n38903, n38904,
         n38905, n38906, n38907, n38908, n38909, n38910, n38911, n38912,
         n38913, n38914, n38915, n38916, n38917, n38918, n38919, n38920;

  DFF_X1 \DRAM_mem_reg[0][31]  ( .D(n9266), .CK(CLK), .Q(n6435), .QN(n37709)
         );
  DFF_X1 \DRAM_mem_reg[0][30]  ( .D(n9265), .CK(CLK), .Q(n6434), .QN(n37708)
         );
  DFF_X1 \DRAM_mem_reg[0][29]  ( .D(n9264), .CK(CLK), .Q(n6433), .QN(n37707)
         );
  DFF_X1 \DRAM_mem_reg[0][28]  ( .D(n9263), .CK(CLK), .Q(n6432), .QN(n37706)
         );
  DFF_X1 \DRAM_mem_reg[0][27]  ( .D(n9262), .CK(CLK), .Q(n6431), .QN(n37705)
         );
  DFF_X1 \DRAM_mem_reg[0][26]  ( .D(n9261), .CK(CLK), .Q(n6430), .QN(n37704)
         );
  DFF_X1 \DRAM_mem_reg[0][25]  ( .D(n9260), .CK(CLK), .Q(n6429), .QN(n37703)
         );
  DFF_X1 \DRAM_mem_reg[0][24]  ( .D(n9259), .CK(CLK), .Q(n6428), .QN(n37702)
         );
  DFF_X1 \DRAM_mem_reg[0][23]  ( .D(n9258), .CK(CLK), .Q(n6427), .QN(n37701)
         );
  DFF_X1 \DRAM_mem_reg[0][22]  ( .D(n9257), .CK(CLK), .Q(n6426), .QN(n37700)
         );
  DFF_X1 \DRAM_mem_reg[0][21]  ( .D(n9256), .CK(CLK), .Q(n6425), .QN(n37699)
         );
  DFF_X1 \DRAM_mem_reg[0][20]  ( .D(n9255), .CK(CLK), .Q(n6424), .QN(n37698)
         );
  DFF_X1 \DRAM_mem_reg[0][19]  ( .D(n9254), .CK(CLK), .Q(n6423), .QN(n37697)
         );
  DFF_X1 \DRAM_mem_reg[0][18]  ( .D(n9253), .CK(CLK), .Q(n6422), .QN(n37696)
         );
  DFF_X1 \DRAM_mem_reg[0][17]  ( .D(n9252), .CK(CLK), .Q(n6421), .QN(n37695)
         );
  DFF_X1 \DRAM_mem_reg[0][16]  ( .D(n9251), .CK(CLK), .Q(n6420), .QN(n37694)
         );
  DFF_X1 \DRAM_mem_reg[0][15]  ( .D(n9250), .CK(CLK), .Q(n6419), .QN(n37693)
         );
  DFF_X1 \DRAM_mem_reg[0][14]  ( .D(n9249), .CK(CLK), .Q(n6418), .QN(n37692)
         );
  DFF_X1 \DRAM_mem_reg[0][13]  ( .D(n9248), .CK(CLK), .Q(n6417), .QN(n37691)
         );
  DFF_X1 \DRAM_mem_reg[0][12]  ( .D(n9247), .CK(CLK), .Q(n6416), .QN(n37690)
         );
  DFF_X1 \DRAM_mem_reg[0][11]  ( .D(n9246), .CK(CLK), .Q(n6415), .QN(n37689)
         );
  DFF_X1 \DRAM_mem_reg[0][10]  ( .D(n9245), .CK(CLK), .Q(n6414), .QN(n37688)
         );
  DFF_X1 \DRAM_mem_reg[0][9]  ( .D(n9244), .CK(CLK), .Q(n6413), .QN(n37687) );
  DFF_X1 \DRAM_mem_reg[0][8]  ( .D(n9243), .CK(CLK), .Q(n6412), .QN(n37686) );
  DFF_X1 \DRAM_mem_reg[0][7]  ( .D(n9242), .CK(CLK), .Q(n6411), .QN(n37685) );
  DFF_X1 \DRAM_mem_reg[0][6]  ( .D(n9241), .CK(CLK), .Q(n6410), .QN(n37684) );
  DFF_X1 \DRAM_mem_reg[0][5]  ( .D(n9240), .CK(CLK), .Q(n6409), .QN(n37683) );
  DFF_X1 \DRAM_mem_reg[0][4]  ( .D(n9239), .CK(CLK), .Q(n6407), .QN(n37682) );
  DFF_X1 \DRAM_mem_reg[0][3]  ( .D(n9238), .CK(CLK), .Q(n6405), .QN(n37681) );
  DFF_X1 \DRAM_mem_reg[0][2]  ( .D(n9237), .CK(CLK), .Q(n6404), .QN(n37680) );
  DFF_X1 \DRAM_mem_reg[0][1]  ( .D(n9236), .CK(CLK), .Q(n6403), .QN(n37679) );
  DFF_X1 \DRAM_mem_reg[0][0]  ( .D(n9235), .CK(CLK), .Q(n6402), .QN(n37678) );
  DFF_X1 \DRAM_mem_reg[1][31]  ( .D(n9234), .CK(CLK), .Q(n5555), .QN(n37549)
         );
  DFF_X1 \DRAM_mem_reg[1][30]  ( .D(n9233), .CK(CLK), .Q(n5606), .QN(n37548)
         );
  DFF_X1 \DRAM_mem_reg[1][29]  ( .D(n9232), .CK(CLK), .Q(n5648), .QN(n37547)
         );
  DFF_X1 \DRAM_mem_reg[1][28]  ( .D(n9231), .CK(CLK), .Q(n5690), .QN(n37546)
         );
  DFF_X1 \DRAM_mem_reg[1][27]  ( .D(n9230), .CK(CLK), .Q(n5732), .QN(n37545)
         );
  DFF_X1 \DRAM_mem_reg[1][26]  ( .D(n9229), .CK(CLK), .Q(n5774), .QN(n37544)
         );
  DFF_X1 \DRAM_mem_reg[1][25]  ( .D(n9228), .CK(CLK), .Q(n5816), .QN(n37543)
         );
  DFF_X1 \DRAM_mem_reg[1][24]  ( .D(n9227), .CK(CLK), .Q(n5858), .QN(n37542)
         );
  DFF_X1 \DRAM_mem_reg[1][23]  ( .D(n9226), .CK(CLK), .Q(n5900), .QN(n37541)
         );
  DFF_X1 \DRAM_mem_reg[1][22]  ( .D(n9225), .CK(CLK), .Q(n5942), .QN(n37540)
         );
  DFF_X1 \DRAM_mem_reg[1][21]  ( .D(n9224), .CK(CLK), .Q(n5984), .QN(n37539)
         );
  DFF_X1 \DRAM_mem_reg[1][20]  ( .D(n9223), .CK(CLK), .Q(n6026), .QN(n37538)
         );
  DFF_X1 \DRAM_mem_reg[1][19]  ( .D(n9222), .CK(CLK), .Q(n6068), .QN(n37537)
         );
  DFF_X1 \DRAM_mem_reg[1][18]  ( .D(n9221), .CK(CLK), .Q(n6110), .QN(n37536)
         );
  DFF_X1 \DRAM_mem_reg[1][17]  ( .D(n9220), .CK(CLK), .Q(n6152), .QN(n37535)
         );
  DFF_X1 \DRAM_mem_reg[1][16]  ( .D(n9219), .CK(CLK), .Q(n6194), .QN(n37534)
         );
  DFF_X1 \DRAM_mem_reg[1][15]  ( .D(n9218), .CK(CLK), .Q(n6236), .QN(n37533)
         );
  DFF_X1 \DRAM_mem_reg[1][14]  ( .D(n9217), .CK(CLK), .Q(n6278), .QN(n37532)
         );
  DFF_X1 \DRAM_mem_reg[1][13]  ( .D(n9216), .CK(CLK), .Q(n6320), .QN(n37531)
         );
  DFF_X1 \DRAM_mem_reg[1][12]  ( .D(n9215), .CK(CLK), .Q(n6362), .QN(n37530)
         );
  DFF_X1 \DRAM_mem_reg[1][11]  ( .D(n9214), .CK(CLK), .Q(n6532), .QN(n37529)
         );
  DFF_X1 \DRAM_mem_reg[1][10]  ( .D(n9213), .CK(CLK), .Q(n6574), .QN(n37528)
         );
  DFF_X1 \DRAM_mem_reg[1][9]  ( .D(n9212), .CK(CLK), .Q(n6616), .QN(n37527) );
  DFF_X1 \DRAM_mem_reg[1][8]  ( .D(n9211), .CK(CLK), .Q(n6658), .QN(n37526) );
  DFF_X1 \DRAM_mem_reg[1][7]  ( .D(n9210), .CK(CLK), .Q(n9292), .QN(n37525) );
  DFF_X1 \DRAM_mem_reg[1][6]  ( .D(n9209), .CK(CLK), .Q(n9334), .QN(n37524) );
  DFF_X1 \DRAM_mem_reg[1][5]  ( .D(n9208), .CK(CLK), .Q(n9376), .QN(n37523) );
  DFF_X1 \DRAM_mem_reg[1][4]  ( .D(n9207), .CK(CLK), .Q(n9418), .QN(n37522) );
  DFF_X1 \DRAM_mem_reg[1][3]  ( .D(n9206), .CK(CLK), .Q(n9460), .QN(n37521) );
  DFF_X1 \DRAM_mem_reg[1][2]  ( .D(n9205), .CK(CLK), .Q(n9502), .QN(n37520) );
  DFF_X1 \DRAM_mem_reg[1][1]  ( .D(n9204), .CK(CLK), .Q(n9544), .QN(n37519) );
  DFF_X1 \DRAM_mem_reg[1][0]  ( .D(n9203), .CK(CLK), .Q(n9605), .QN(n37518) );
  DFF_X1 \DRAM_mem_reg[2][31]  ( .D(n9202), .CK(CLK), .QN(n35709) );
  DFF_X1 \DRAM_mem_reg[2][30]  ( .D(n9201), .CK(CLK), .QN(n35708) );
  DFF_X1 \DRAM_mem_reg[2][29]  ( .D(n9200), .CK(CLK), .QN(n35707) );
  DFF_X1 \DRAM_mem_reg[2][28]  ( .D(n9199), .CK(CLK), .QN(n35706) );
  DFF_X1 \DRAM_mem_reg[2][27]  ( .D(n9198), .CK(CLK), .QN(n35705) );
  DFF_X1 \DRAM_mem_reg[2][26]  ( .D(n9197), .CK(CLK), .QN(n35704) );
  DFF_X1 \DRAM_mem_reg[2][25]  ( .D(n9196), .CK(CLK), .QN(n35703) );
  DFF_X1 \DRAM_mem_reg[2][24]  ( .D(n9195), .CK(CLK), .QN(n35702) );
  DFF_X1 \DRAM_mem_reg[2][23]  ( .D(n9194), .CK(CLK), .QN(n35853) );
  DFF_X1 \DRAM_mem_reg[2][22]  ( .D(n9193), .CK(CLK), .QN(n35852) );
  DFF_X1 \DRAM_mem_reg[2][21]  ( .D(n9192), .CK(CLK), .QN(n35851) );
  DFF_X1 \DRAM_mem_reg[2][20]  ( .D(n9191), .CK(CLK), .QN(n35850) );
  DFF_X1 \DRAM_mem_reg[2][19]  ( .D(n9190), .CK(CLK), .QN(n35849) );
  DFF_X1 \DRAM_mem_reg[2][18]  ( .D(n9189), .CK(CLK), .QN(n35848) );
  DFF_X1 \DRAM_mem_reg[2][17]  ( .D(n9188), .CK(CLK), .QN(n35847) );
  DFF_X1 \DRAM_mem_reg[2][16]  ( .D(n9187), .CK(CLK), .QN(n35846) );
  DFF_X1 \DRAM_mem_reg[2][15]  ( .D(n9186), .CK(CLK), .QN(n35845) );
  DFF_X1 \DRAM_mem_reg[2][14]  ( .D(n9185), .CK(CLK), .QN(n35844) );
  DFF_X1 \DRAM_mem_reg[2][13]  ( .D(n9184), .CK(CLK), .QN(n35843) );
  DFF_X1 \DRAM_mem_reg[2][12]  ( .D(n9183), .CK(CLK), .QN(n35842) );
  DFF_X1 \DRAM_mem_reg[2][11]  ( .D(n9182), .CK(CLK), .QN(n35841) );
  DFF_X1 \DRAM_mem_reg[2][10]  ( .D(n9181), .CK(CLK), .QN(n35840) );
  DFF_X1 \DRAM_mem_reg[2][9]  ( .D(n9180), .CK(CLK), .QN(n35839) );
  DFF_X1 \DRAM_mem_reg[2][8]  ( .D(n9179), .CK(CLK), .QN(n35838) );
  DFF_X1 \DRAM_mem_reg[2][7]  ( .D(n9178), .CK(CLK), .QN(n35837) );
  DFF_X1 \DRAM_mem_reg[2][6]  ( .D(n9177), .CK(CLK), .QN(n35836) );
  DFF_X1 \DRAM_mem_reg[2][5]  ( .D(n9176), .CK(CLK), .QN(n35835) );
  DFF_X1 \DRAM_mem_reg[2][4]  ( .D(n9175), .CK(CLK), .QN(n35834) );
  DFF_X1 \DRAM_mem_reg[2][3]  ( .D(n9174), .CK(CLK), .QN(n35833) );
  DFF_X1 \DRAM_mem_reg[2][2]  ( .D(n9173), .CK(CLK), .QN(n35832) );
  DFF_X1 \DRAM_mem_reg[2][1]  ( .D(n9172), .CK(CLK), .QN(n35831) );
  DFF_X1 \DRAM_mem_reg[2][0]  ( .D(n9171), .CK(CLK), .QN(n35830) );
  DFF_X1 \DRAM_mem_reg[3][31]  ( .D(n9170), .CK(CLK), .QN(n36221) );
  DFF_X1 \DRAM_mem_reg[3][30]  ( .D(n9169), .CK(CLK), .QN(n36220) );
  DFF_X1 \DRAM_mem_reg[3][29]  ( .D(n9168), .CK(CLK), .QN(n36219) );
  DFF_X1 \DRAM_mem_reg[3][28]  ( .D(n9167), .CK(CLK), .QN(n36218) );
  DFF_X1 \DRAM_mem_reg[3][27]  ( .D(n9166), .CK(CLK), .QN(n36217) );
  DFF_X1 \DRAM_mem_reg[3][26]  ( .D(n9165), .CK(CLK), .QN(n36216) );
  DFF_X1 \DRAM_mem_reg[3][25]  ( .D(n9164), .CK(CLK), .QN(n36215) );
  DFF_X1 \DRAM_mem_reg[3][24]  ( .D(n9163), .CK(CLK), .QN(n36214) );
  DFF_X1 \DRAM_mem_reg[3][23]  ( .D(n9162), .CK(CLK), .QN(n36365) );
  DFF_X1 \DRAM_mem_reg[3][22]  ( .D(n9161), .CK(CLK), .QN(n36364) );
  DFF_X1 \DRAM_mem_reg[3][21]  ( .D(n9160), .CK(CLK), .QN(n36363) );
  DFF_X1 \DRAM_mem_reg[3][20]  ( .D(n9159), .CK(CLK), .QN(n36362) );
  DFF_X1 \DRAM_mem_reg[3][19]  ( .D(n9158), .CK(CLK), .QN(n36361) );
  DFF_X1 \DRAM_mem_reg[3][18]  ( .D(n9157), .CK(CLK), .QN(n36360) );
  DFF_X1 \DRAM_mem_reg[3][17]  ( .D(n9156), .CK(CLK), .QN(n36359) );
  DFF_X1 \DRAM_mem_reg[3][16]  ( .D(n9155), .CK(CLK), .QN(n36358) );
  DFF_X1 \DRAM_mem_reg[3][15]  ( .D(n9154), .CK(CLK), .QN(n36357) );
  DFF_X1 \DRAM_mem_reg[3][14]  ( .D(n9153), .CK(CLK), .QN(n36356) );
  DFF_X1 \DRAM_mem_reg[3][13]  ( .D(n9152), .CK(CLK), .QN(n36355) );
  DFF_X1 \DRAM_mem_reg[3][12]  ( .D(n9151), .CK(CLK), .QN(n36354) );
  DFF_X1 \DRAM_mem_reg[3][11]  ( .D(n9150), .CK(CLK), .QN(n36353) );
  DFF_X1 \DRAM_mem_reg[3][10]  ( .D(n9149), .CK(CLK), .QN(n36352) );
  DFF_X1 \DRAM_mem_reg[3][9]  ( .D(n9148), .CK(CLK), .QN(n36351) );
  DFF_X1 \DRAM_mem_reg[3][8]  ( .D(n9147), .CK(CLK), .QN(n36350) );
  DFF_X1 \DRAM_mem_reg[3][7]  ( .D(n9146), .CK(CLK), .QN(n36349) );
  DFF_X1 \DRAM_mem_reg[3][6]  ( .D(n9145), .CK(CLK), .QN(n36348) );
  DFF_X1 \DRAM_mem_reg[3][5]  ( .D(n9144), .CK(CLK), .QN(n36347) );
  DFF_X1 \DRAM_mem_reg[3][4]  ( .D(n9143), .CK(CLK), .QN(n36346) );
  DFF_X1 \DRAM_mem_reg[3][3]  ( .D(n9142), .CK(CLK), .QN(n36345) );
  DFF_X1 \DRAM_mem_reg[3][2]  ( .D(n9141), .CK(CLK), .QN(n36344) );
  DFF_X1 \DRAM_mem_reg[3][1]  ( .D(n9140), .CK(CLK), .QN(n36343) );
  DFF_X1 \DRAM_mem_reg[3][0]  ( .D(n9139), .CK(CLK), .QN(n36342) );
  DFF_X1 \DRAM_mem_reg[4][31]  ( .D(n9138), .CK(CLK), .QN(n35197) );
  DFF_X1 \DRAM_mem_reg[4][30]  ( .D(n9137), .CK(CLK), .QN(n35196) );
  DFF_X1 \DRAM_mem_reg[4][29]  ( .D(n9136), .CK(CLK), .QN(n35195) );
  DFF_X1 \DRAM_mem_reg[4][28]  ( .D(n9135), .CK(CLK), .QN(n35194) );
  DFF_X1 \DRAM_mem_reg[4][27]  ( .D(n9134), .CK(CLK), .QN(n35193) );
  DFF_X1 \DRAM_mem_reg[4][26]  ( .D(n9133), .CK(CLK), .QN(n35192) );
  DFF_X1 \DRAM_mem_reg[4][25]  ( .D(n9132), .CK(CLK), .QN(n35191) );
  DFF_X1 \DRAM_mem_reg[4][24]  ( .D(n9131), .CK(CLK), .QN(n35190) );
  DFF_X1 \DRAM_mem_reg[4][23]  ( .D(n9130), .CK(CLK), .QN(n35341) );
  DFF_X1 \DRAM_mem_reg[4][22]  ( .D(n9129), .CK(CLK), .QN(n35340) );
  DFF_X1 \DRAM_mem_reg[4][21]  ( .D(n9128), .CK(CLK), .QN(n35339) );
  DFF_X1 \DRAM_mem_reg[4][20]  ( .D(n9127), .CK(CLK), .QN(n35338) );
  DFF_X1 \DRAM_mem_reg[4][19]  ( .D(n9126), .CK(CLK), .QN(n35337) );
  DFF_X1 \DRAM_mem_reg[4][18]  ( .D(n9125), .CK(CLK), .QN(n35336) );
  DFF_X1 \DRAM_mem_reg[4][17]  ( .D(n9124), .CK(CLK), .QN(n35335) );
  DFF_X1 \DRAM_mem_reg[4][16]  ( .D(n9123), .CK(CLK), .QN(n35334) );
  DFF_X1 \DRAM_mem_reg[4][15]  ( .D(n9122), .CK(CLK), .QN(n35333) );
  DFF_X1 \DRAM_mem_reg[4][14]  ( .D(n9121), .CK(CLK), .QN(n35332) );
  DFF_X1 \DRAM_mem_reg[4][13]  ( .D(n9120), .CK(CLK), .QN(n35331) );
  DFF_X1 \DRAM_mem_reg[4][12]  ( .D(n9119), .CK(CLK), .QN(n35330) );
  DFF_X1 \DRAM_mem_reg[4][11]  ( .D(n9118), .CK(CLK), .QN(n35329) );
  DFF_X1 \DRAM_mem_reg[4][10]  ( .D(n9117), .CK(CLK), .QN(n35328) );
  DFF_X1 \DRAM_mem_reg[4][9]  ( .D(n9116), .CK(CLK), .QN(n35327) );
  DFF_X1 \DRAM_mem_reg[4][8]  ( .D(n9115), .CK(CLK), .QN(n35326) );
  DFF_X1 \DRAM_mem_reg[4][7]  ( .D(n9114), .CK(CLK), .QN(n35325) );
  DFF_X1 \DRAM_mem_reg[4][6]  ( .D(n9113), .CK(CLK), .QN(n35324) );
  DFF_X1 \DRAM_mem_reg[4][5]  ( .D(n9112), .CK(CLK), .QN(n35323) );
  DFF_X1 \DRAM_mem_reg[4][4]  ( .D(n9111), .CK(CLK), .QN(n35322) );
  DFF_X1 \DRAM_mem_reg[4][3]  ( .D(n9110), .CK(CLK), .QN(n35321) );
  DFF_X1 \DRAM_mem_reg[4][2]  ( .D(n9109), .CK(CLK), .QN(n35320) );
  DFF_X1 \DRAM_mem_reg[4][1]  ( .D(n9108), .CK(CLK), .QN(n35319) );
  DFF_X1 \DRAM_mem_reg[4][0]  ( .D(n9107), .CK(CLK), .QN(n35318) );
  DFF_X1 \DRAM_mem_reg[5][31]  ( .D(n9106), .CK(CLK), .Q(n6401), .QN(n37677)
         );
  DFF_X1 \DRAM_mem_reg[5][30]  ( .D(n9105), .CK(CLK), .Q(n6400), .QN(n37676)
         );
  DFF_X1 \DRAM_mem_reg[5][29]  ( .D(n9104), .CK(CLK), .Q(n6399), .QN(n37675)
         );
  DFF_X1 \DRAM_mem_reg[5][28]  ( .D(n9103), .CK(CLK), .Q(n6398), .QN(n37674)
         );
  DFF_X1 \DRAM_mem_reg[5][27]  ( .D(n9102), .CK(CLK), .Q(n6397), .QN(n37673)
         );
  DFF_X1 \DRAM_mem_reg[5][26]  ( .D(n9101), .CK(CLK), .Q(n6396), .QN(n37672)
         );
  DFF_X1 \DRAM_mem_reg[5][25]  ( .D(n9100), .CK(CLK), .Q(n6395), .QN(n37671)
         );
  DFF_X1 \DRAM_mem_reg[5][24]  ( .D(n9099), .CK(CLK), .Q(n6394), .QN(n37670)
         );
  DFF_X1 \DRAM_mem_reg[5][23]  ( .D(n9098), .CK(CLK), .Q(n6393), .QN(n37669)
         );
  DFF_X1 \DRAM_mem_reg[5][22]  ( .D(n9097), .CK(CLK), .Q(n6392), .QN(n37668)
         );
  DFF_X1 \DRAM_mem_reg[5][21]  ( .D(n9096), .CK(CLK), .Q(n6391), .QN(n37667)
         );
  DFF_X1 \DRAM_mem_reg[5][20]  ( .D(n9095), .CK(CLK), .Q(n6390), .QN(n37666)
         );
  DFF_X1 \DRAM_mem_reg[5][19]  ( .D(n9094), .CK(CLK), .Q(n6389), .QN(n37665)
         );
  DFF_X1 \DRAM_mem_reg[5][18]  ( .D(n9093), .CK(CLK), .Q(n6388), .QN(n37664)
         );
  DFF_X1 \DRAM_mem_reg[5][17]  ( .D(n9092), .CK(CLK), .Q(n6387), .QN(n37663)
         );
  DFF_X1 \DRAM_mem_reg[5][16]  ( .D(n9091), .CK(CLK), .Q(n6386), .QN(n37662)
         );
  DFF_X1 \DRAM_mem_reg[5][15]  ( .D(n9090), .CK(CLK), .Q(n6385), .QN(n37661)
         );
  DFF_X1 \DRAM_mem_reg[5][14]  ( .D(n9089), .CK(CLK), .Q(n6384), .QN(n37660)
         );
  DFF_X1 \DRAM_mem_reg[5][13]  ( .D(n9088), .CK(CLK), .Q(n6383), .QN(n37659)
         );
  DFF_X1 \DRAM_mem_reg[5][12]  ( .D(n9087), .CK(CLK), .Q(n6382), .QN(n37658)
         );
  DFF_X1 \DRAM_mem_reg[5][11]  ( .D(n9086), .CK(CLK), .Q(n6381), .QN(n37657)
         );
  DFF_X1 \DRAM_mem_reg[5][10]  ( .D(n9085), .CK(CLK), .Q(n6380), .QN(n37656)
         );
  DFF_X1 \DRAM_mem_reg[5][9]  ( .D(n9084), .CK(CLK), .Q(n6379), .QN(n37655) );
  DFF_X1 \DRAM_mem_reg[5][8]  ( .D(n9083), .CK(CLK), .Q(n6378), .QN(n37654) );
  DFF_X1 \DRAM_mem_reg[5][7]  ( .D(n9082), .CK(CLK), .Q(n6377), .QN(n37653) );
  DFF_X1 \DRAM_mem_reg[5][6]  ( .D(n9081), .CK(CLK), .Q(n6376), .QN(n37652) );
  DFF_X1 \DRAM_mem_reg[5][5]  ( .D(n9080), .CK(CLK), .Q(n6375), .QN(n37651) );
  DFF_X1 \DRAM_mem_reg[5][4]  ( .D(n9079), .CK(CLK), .Q(n6374), .QN(n37650) );
  DFF_X1 \DRAM_mem_reg[5][3]  ( .D(n9078), .CK(CLK), .Q(n6372), .QN(n37649) );
  DFF_X1 \DRAM_mem_reg[5][2]  ( .D(n9077), .CK(CLK), .Q(n6370), .QN(n37648) );
  DFF_X1 \DRAM_mem_reg[5][1]  ( .D(n9076), .CK(CLK), .Q(n6369), .QN(n37647) );
  DFF_X1 \DRAM_mem_reg[5][0]  ( .D(n9075), .CK(CLK), .Q(n6368), .QN(n37646) );
  DFF_X1 \DRAM_mem_reg[6][31]  ( .D(n9074), .CK(CLK), .Q(n5553), .QN(n37517)
         );
  DFF_X1 \DRAM_mem_reg[6][30]  ( .D(n9073), .CK(CLK), .Q(n5604), .QN(n37516)
         );
  DFF_X1 \DRAM_mem_reg[6][29]  ( .D(n9072), .CK(CLK), .Q(n5646), .QN(n37515)
         );
  DFF_X1 \DRAM_mem_reg[6][28]  ( .D(n9071), .CK(CLK), .Q(n5688), .QN(n37514)
         );
  DFF_X1 \DRAM_mem_reg[6][27]  ( .D(n9070), .CK(CLK), .Q(n5730), .QN(n37513)
         );
  DFF_X1 \DRAM_mem_reg[6][26]  ( .D(n9069), .CK(CLK), .Q(n5772), .QN(n37512)
         );
  DFF_X1 \DRAM_mem_reg[6][25]  ( .D(n9068), .CK(CLK), .Q(n5814), .QN(n37511)
         );
  DFF_X1 \DRAM_mem_reg[6][24]  ( .D(n9067), .CK(CLK), .Q(n5856), .QN(n37510)
         );
  DFF_X1 \DRAM_mem_reg[6][23]  ( .D(n9066), .CK(CLK), .Q(n5898), .QN(n37509)
         );
  DFF_X1 \DRAM_mem_reg[6][22]  ( .D(n9065), .CK(CLK), .Q(n5940), .QN(n37508)
         );
  DFF_X1 \DRAM_mem_reg[6][21]  ( .D(n9064), .CK(CLK), .Q(n5982), .QN(n37507)
         );
  DFF_X1 \DRAM_mem_reg[6][20]  ( .D(n9063), .CK(CLK), .Q(n6024), .QN(n37506)
         );
  DFF_X1 \DRAM_mem_reg[6][19]  ( .D(n9062), .CK(CLK), .Q(n6066), .QN(n37505)
         );
  DFF_X1 \DRAM_mem_reg[6][18]  ( .D(n9061), .CK(CLK), .Q(n6108), .QN(n37504)
         );
  DFF_X1 \DRAM_mem_reg[6][17]  ( .D(n9060), .CK(CLK), .Q(n6150), .QN(n37503)
         );
  DFF_X1 \DRAM_mem_reg[6][16]  ( .D(n9059), .CK(CLK), .Q(n6192), .QN(n37502)
         );
  DFF_X1 \DRAM_mem_reg[6][15]  ( .D(n9058), .CK(CLK), .Q(n6234), .QN(n37501)
         );
  DFF_X1 \DRAM_mem_reg[6][14]  ( .D(n9057), .CK(CLK), .Q(n6276), .QN(n37500)
         );
  DFF_X1 \DRAM_mem_reg[6][13]  ( .D(n9056), .CK(CLK), .Q(n6318), .QN(n37499)
         );
  DFF_X1 \DRAM_mem_reg[6][12]  ( .D(n9055), .CK(CLK), .Q(n6360), .QN(n37498)
         );
  DFF_X1 \DRAM_mem_reg[6][11]  ( .D(n9054), .CK(CLK), .Q(n6530), .QN(n37497)
         );
  DFF_X1 \DRAM_mem_reg[6][10]  ( .D(n9053), .CK(CLK), .Q(n6572), .QN(n37496)
         );
  DFF_X1 \DRAM_mem_reg[6][9]  ( .D(n9052), .CK(CLK), .Q(n6614), .QN(n37495) );
  DFF_X1 \DRAM_mem_reg[6][8]  ( .D(n9051), .CK(CLK), .Q(n6656), .QN(n37494) );
  DFF_X1 \DRAM_mem_reg[6][7]  ( .D(n9050), .CK(CLK), .Q(n9290), .QN(n37493) );
  DFF_X1 \DRAM_mem_reg[6][6]  ( .D(n9049), .CK(CLK), .Q(n9332), .QN(n37492) );
  DFF_X1 \DRAM_mem_reg[6][5]  ( .D(n9048), .CK(CLK), .Q(n9374), .QN(n37491) );
  DFF_X1 \DRAM_mem_reg[6][4]  ( .D(n9047), .CK(CLK), .Q(n9416), .QN(n37490) );
  DFF_X1 \DRAM_mem_reg[6][3]  ( .D(n9046), .CK(CLK), .Q(n9458), .QN(n37489) );
  DFF_X1 \DRAM_mem_reg[6][2]  ( .D(n9045), .CK(CLK), .Q(n9500), .QN(n37488) );
  DFF_X1 \DRAM_mem_reg[6][1]  ( .D(n9044), .CK(CLK), .Q(n9542), .QN(n37487) );
  DFF_X1 \DRAM_mem_reg[6][0]  ( .D(n9043), .CK(CLK), .Q(n9602), .QN(n37486) );
  DFF_X1 \DRAM_mem_reg[7][31]  ( .D(n9042), .CK(CLK), .QN(n36029) );
  DFF_X1 \DRAM_mem_reg[7][30]  ( .D(n9041), .CK(CLK), .QN(n36028) );
  DFF_X1 \DRAM_mem_reg[7][29]  ( .D(n9040), .CK(CLK), .QN(n36027) );
  DFF_X1 \DRAM_mem_reg[7][28]  ( .D(n9039), .CK(CLK), .QN(n36026) );
  DFF_X1 \DRAM_mem_reg[7][27]  ( .D(n9038), .CK(CLK), .QN(n36025) );
  DFF_X1 \DRAM_mem_reg[7][26]  ( .D(n9037), .CK(CLK), .QN(n36024) );
  DFF_X1 \DRAM_mem_reg[7][25]  ( .D(n9036), .CK(CLK), .QN(n36023) );
  DFF_X1 \DRAM_mem_reg[7][24]  ( .D(n9035), .CK(CLK), .QN(n36022) );
  DFF_X1 \DRAM_mem_reg[7][23]  ( .D(n9034), .CK(CLK), .QN(n36019) );
  DFF_X1 \DRAM_mem_reg[7][22]  ( .D(n9033), .CK(CLK), .QN(n36015) );
  DFF_X1 \DRAM_mem_reg[7][21]  ( .D(n9032), .CK(CLK), .QN(n36011) );
  DFF_X1 \DRAM_mem_reg[7][20]  ( .D(n9031), .CK(CLK), .QN(n36007) );
  DFF_X1 \DRAM_mem_reg[7][19]  ( .D(n9030), .CK(CLK), .QN(n36003) );
  DFF_X1 \DRAM_mem_reg[7][18]  ( .D(n9029), .CK(CLK), .QN(n35999) );
  DFF_X1 \DRAM_mem_reg[7][17]  ( .D(n9028), .CK(CLK), .QN(n35995) );
  DFF_X1 \DRAM_mem_reg[7][16]  ( .D(n9027), .CK(CLK), .QN(n35991) );
  DFF_X1 \DRAM_mem_reg[7][15]  ( .D(n9026), .CK(CLK), .QN(n35987) );
  DFF_X1 \DRAM_mem_reg[7][14]  ( .D(n9025), .CK(CLK), .QN(n35983) );
  DFF_X1 \DRAM_mem_reg[7][13]  ( .D(n9024), .CK(CLK), .QN(n35979) );
  DFF_X1 \DRAM_mem_reg[7][12]  ( .D(n9023), .CK(CLK), .QN(n35975) );
  DFF_X1 \DRAM_mem_reg[7][11]  ( .D(n9022), .CK(CLK), .QN(n35971) );
  DFF_X1 \DRAM_mem_reg[7][10]  ( .D(n9021), .CK(CLK), .QN(n35967) );
  DFF_X1 \DRAM_mem_reg[7][9]  ( .D(n9020), .CK(CLK), .QN(n35963) );
  DFF_X1 \DRAM_mem_reg[7][8]  ( .D(n9019), .CK(CLK), .QN(n35959) );
  DFF_X1 \DRAM_mem_reg[7][7]  ( .D(n9018), .CK(CLK), .QN(n35955) );
  DFF_X1 \DRAM_mem_reg[7][6]  ( .D(n9017), .CK(CLK), .QN(n35951) );
  DFF_X1 \DRAM_mem_reg[7][5]  ( .D(n9016), .CK(CLK), .QN(n35947) );
  DFF_X1 \DRAM_mem_reg[7][4]  ( .D(n9015), .CK(CLK), .QN(n35943) );
  DFF_X1 \DRAM_mem_reg[7][3]  ( .D(n9014), .CK(CLK), .QN(n35939) );
  DFF_X1 \DRAM_mem_reg[7][2]  ( .D(n9013), .CK(CLK), .QN(n35935) );
  DFF_X1 \DRAM_mem_reg[7][1]  ( .D(n9012), .CK(CLK), .QN(n35931) );
  DFF_X1 \DRAM_mem_reg[7][0]  ( .D(n9011), .CK(CLK), .QN(n35927) );
  DFF_X1 \DRAM_mem_reg[8][31]  ( .D(n9010), .CK(CLK), .QN(n36541) );
  DFF_X1 \DRAM_mem_reg[8][30]  ( .D(n9009), .CK(CLK), .QN(n36540) );
  DFF_X1 \DRAM_mem_reg[8][29]  ( .D(n9008), .CK(CLK), .QN(n36539) );
  DFF_X1 \DRAM_mem_reg[8][28]  ( .D(n9007), .CK(CLK), .QN(n36538) );
  DFF_X1 \DRAM_mem_reg[8][27]  ( .D(n9006), .CK(CLK), .QN(n36537) );
  DFF_X1 \DRAM_mem_reg[8][26]  ( .D(n9005), .CK(CLK), .QN(n36536) );
  DFF_X1 \DRAM_mem_reg[8][25]  ( .D(n9004), .CK(CLK), .QN(n36535) );
  DFF_X1 \DRAM_mem_reg[8][24]  ( .D(n9003), .CK(CLK), .QN(n36534) );
  DFF_X1 \DRAM_mem_reg[8][23]  ( .D(n9002), .CK(CLK), .QN(n36531) );
  DFF_X1 \DRAM_mem_reg[8][22]  ( .D(n9001), .CK(CLK), .QN(n36527) );
  DFF_X1 \DRAM_mem_reg[8][21]  ( .D(n9000), .CK(CLK), .QN(n36523) );
  DFF_X1 \DRAM_mem_reg[8][20]  ( .D(n8999), .CK(CLK), .QN(n36519) );
  DFF_X1 \DRAM_mem_reg[8][19]  ( .D(n8998), .CK(CLK), .QN(n36515) );
  DFF_X1 \DRAM_mem_reg[8][18]  ( .D(n8997), .CK(CLK), .QN(n36511) );
  DFF_X1 \DRAM_mem_reg[8][17]  ( .D(n8996), .CK(CLK), .QN(n36507) );
  DFF_X1 \DRAM_mem_reg[8][16]  ( .D(n8995), .CK(CLK), .QN(n36503) );
  DFF_X1 \DRAM_mem_reg[8][15]  ( .D(n8994), .CK(CLK), .QN(n36499) );
  DFF_X1 \DRAM_mem_reg[8][14]  ( .D(n8993), .CK(CLK), .QN(n36495) );
  DFF_X1 \DRAM_mem_reg[8][13]  ( .D(n8992), .CK(CLK), .QN(n36491) );
  DFF_X1 \DRAM_mem_reg[8][12]  ( .D(n8991), .CK(CLK), .QN(n36487) );
  DFF_X1 \DRAM_mem_reg[8][11]  ( .D(n8990), .CK(CLK), .QN(n36483) );
  DFF_X1 \DRAM_mem_reg[8][10]  ( .D(n8989), .CK(CLK), .QN(n36479) );
  DFF_X1 \DRAM_mem_reg[8][9]  ( .D(n8988), .CK(CLK), .QN(n36475) );
  DFF_X1 \DRAM_mem_reg[8][8]  ( .D(n8987), .CK(CLK), .QN(n36471) );
  DFF_X1 \DRAM_mem_reg[8][7]  ( .D(n8986), .CK(CLK), .QN(n36467) );
  DFF_X1 \DRAM_mem_reg[8][6]  ( .D(n8985), .CK(CLK), .QN(n36463) );
  DFF_X1 \DRAM_mem_reg[8][5]  ( .D(n8984), .CK(CLK), .QN(n36459) );
  DFF_X1 \DRAM_mem_reg[8][4]  ( .D(n8983), .CK(CLK), .QN(n36455) );
  DFF_X1 \DRAM_mem_reg[8][3]  ( .D(n8982), .CK(CLK), .QN(n36451) );
  DFF_X1 \DRAM_mem_reg[8][2]  ( .D(n8981), .CK(CLK), .QN(n36447) );
  DFF_X1 \DRAM_mem_reg[8][1]  ( .D(n8980), .CK(CLK), .QN(n36443) );
  DFF_X1 \DRAM_mem_reg[8][0]  ( .D(n8979), .CK(CLK), .QN(n36439) );
  DFF_X1 \DRAM_mem_reg[9][31]  ( .D(n8978), .CK(CLK), .QN(n35517) );
  DFF_X1 \DRAM_mem_reg[9][30]  ( .D(n8977), .CK(CLK), .QN(n35516) );
  DFF_X1 \DRAM_mem_reg[9][29]  ( .D(n8976), .CK(CLK), .QN(n35515) );
  DFF_X1 \DRAM_mem_reg[9][28]  ( .D(n8975), .CK(CLK), .QN(n35514) );
  DFF_X1 \DRAM_mem_reg[9][27]  ( .D(n8974), .CK(CLK), .QN(n35513) );
  DFF_X1 \DRAM_mem_reg[9][26]  ( .D(n8973), .CK(CLK), .QN(n35512) );
  DFF_X1 \DRAM_mem_reg[9][25]  ( .D(n8972), .CK(CLK), .QN(n35511) );
  DFF_X1 \DRAM_mem_reg[9][24]  ( .D(n8971), .CK(CLK), .QN(n35510) );
  DFF_X1 \DRAM_mem_reg[9][23]  ( .D(n8970), .CK(CLK), .QN(n35507) );
  DFF_X1 \DRAM_mem_reg[9][22]  ( .D(n8969), .CK(CLK), .QN(n35503) );
  DFF_X1 \DRAM_mem_reg[9][21]  ( .D(n8968), .CK(CLK), .QN(n35499) );
  DFF_X1 \DRAM_mem_reg[9][20]  ( .D(n8967), .CK(CLK), .QN(n35495) );
  DFF_X1 \DRAM_mem_reg[9][19]  ( .D(n8966), .CK(CLK), .QN(n35491) );
  DFF_X1 \DRAM_mem_reg[9][18]  ( .D(n8965), .CK(CLK), .QN(n35487) );
  DFF_X1 \DRAM_mem_reg[9][17]  ( .D(n8964), .CK(CLK), .QN(n35483) );
  DFF_X1 \DRAM_mem_reg[9][16]  ( .D(n8963), .CK(CLK), .QN(n35479) );
  DFF_X1 \DRAM_mem_reg[9][15]  ( .D(n8962), .CK(CLK), .QN(n35475) );
  DFF_X1 \DRAM_mem_reg[9][14]  ( .D(n8961), .CK(CLK), .QN(n35471) );
  DFF_X1 \DRAM_mem_reg[9][13]  ( .D(n8960), .CK(CLK), .QN(n35467) );
  DFF_X1 \DRAM_mem_reg[9][12]  ( .D(n8959), .CK(CLK), .QN(n35463) );
  DFF_X1 \DRAM_mem_reg[9][11]  ( .D(n8958), .CK(CLK), .QN(n35459) );
  DFF_X1 \DRAM_mem_reg[9][10]  ( .D(n8957), .CK(CLK), .QN(n35455) );
  DFF_X1 \DRAM_mem_reg[9][9]  ( .D(n8956), .CK(CLK), .QN(n35451) );
  DFF_X1 \DRAM_mem_reg[9][8]  ( .D(n8955), .CK(CLK), .QN(n35447) );
  DFF_X1 \DRAM_mem_reg[9][7]  ( .D(n8954), .CK(CLK), .QN(n35443) );
  DFF_X1 \DRAM_mem_reg[9][6]  ( .D(n8953), .CK(CLK), .QN(n35439) );
  DFF_X1 \DRAM_mem_reg[9][5]  ( .D(n8952), .CK(CLK), .QN(n35435) );
  DFF_X1 \DRAM_mem_reg[9][4]  ( .D(n8951), .CK(CLK), .QN(n35431) );
  DFF_X1 \DRAM_mem_reg[9][3]  ( .D(n8950), .CK(CLK), .QN(n35427) );
  DFF_X1 \DRAM_mem_reg[9][2]  ( .D(n8949), .CK(CLK), .QN(n35423) );
  DFF_X1 \DRAM_mem_reg[9][1]  ( .D(n8948), .CK(CLK), .QN(n35419) );
  DFF_X1 \DRAM_mem_reg[9][0]  ( .D(n8947), .CK(CLK), .QN(n35415) );
  DFF_X1 \DRAM_mem_reg[10][31]  ( .D(n8946), .CK(CLK), .Q(n6507), .QN(n37645)
         );
  DFF_X1 \DRAM_mem_reg[10][30]  ( .D(n8945), .CK(CLK), .Q(n6506), .QN(n37644)
         );
  DFF_X1 \DRAM_mem_reg[10][29]  ( .D(n8944), .CK(CLK), .Q(n6505), .QN(n37643)
         );
  DFF_X1 \DRAM_mem_reg[10][28]  ( .D(n8943), .CK(CLK), .Q(n6504), .QN(n37642)
         );
  DFF_X1 \DRAM_mem_reg[10][27]  ( .D(n8942), .CK(CLK), .Q(n6503), .QN(n37641)
         );
  DFF_X1 \DRAM_mem_reg[10][26]  ( .D(n8941), .CK(CLK), .Q(n6502), .QN(n37640)
         );
  DFF_X1 \DRAM_mem_reg[10][25]  ( .D(n8940), .CK(CLK), .Q(n6501), .QN(n37639)
         );
  DFF_X1 \DRAM_mem_reg[10][24]  ( .D(n8939), .CK(CLK), .Q(n6500), .QN(n37638)
         );
  DFF_X1 \DRAM_mem_reg[10][23]  ( .D(n8938), .CK(CLK), .Q(n6499), .QN(n37637)
         );
  DFF_X1 \DRAM_mem_reg[10][22]  ( .D(n8937), .CK(CLK), .Q(n6498), .QN(n37636)
         );
  DFF_X1 \DRAM_mem_reg[10][21]  ( .D(n8936), .CK(CLK), .Q(n6497), .QN(n37635)
         );
  DFF_X1 \DRAM_mem_reg[10][20]  ( .D(n8935), .CK(CLK), .Q(n6496), .QN(n37634)
         );
  DFF_X1 \DRAM_mem_reg[10][19]  ( .D(n8934), .CK(CLK), .Q(n6495), .QN(n37633)
         );
  DFF_X1 \DRAM_mem_reg[10][18]  ( .D(n8933), .CK(CLK), .Q(n6494), .QN(n37632)
         );
  DFF_X1 \DRAM_mem_reg[10][17]  ( .D(n8932), .CK(CLK), .Q(n6493), .QN(n37631)
         );
  DFF_X1 \DRAM_mem_reg[10][16]  ( .D(n8931), .CK(CLK), .Q(n6492), .QN(n37630)
         );
  DFF_X1 \DRAM_mem_reg[10][15]  ( .D(n8930), .CK(CLK), .Q(n6491), .QN(n37629)
         );
  DFF_X1 \DRAM_mem_reg[10][14]  ( .D(n8929), .CK(CLK), .Q(n6490), .QN(n37628)
         );
  DFF_X1 \DRAM_mem_reg[10][13]  ( .D(n8928), .CK(CLK), .Q(n6489), .QN(n37627)
         );
  DFF_X1 \DRAM_mem_reg[10][12]  ( .D(n8927), .CK(CLK), .Q(n6488), .QN(n37626)
         );
  DFF_X1 \DRAM_mem_reg[10][11]  ( .D(n8926), .CK(CLK), .Q(n6487), .QN(n37625)
         );
  DFF_X1 \DRAM_mem_reg[10][10]  ( .D(n8925), .CK(CLK), .Q(n6486), .QN(n37624)
         );
  DFF_X1 \DRAM_mem_reg[10][9]  ( .D(n8924), .CK(CLK), .Q(n6485), .QN(n37623)
         );
  DFF_X1 \DRAM_mem_reg[10][8]  ( .D(n8923), .CK(CLK), .Q(n6483), .QN(n37622)
         );
  DFF_X1 \DRAM_mem_reg[10][7]  ( .D(n8922), .CK(CLK), .Q(n6481), .QN(n37621)
         );
  DFF_X1 \DRAM_mem_reg[10][6]  ( .D(n8921), .CK(CLK), .Q(n6480), .QN(n37620)
         );
  DFF_X1 \DRAM_mem_reg[10][5]  ( .D(n8920), .CK(CLK), .Q(n6479), .QN(n37619)
         );
  DFF_X1 \DRAM_mem_reg[10][4]  ( .D(n8919), .CK(CLK), .Q(n6478), .QN(n37618)
         );
  DFF_X1 \DRAM_mem_reg[10][3]  ( .D(n8918), .CK(CLK), .Q(n6477), .QN(n37617)
         );
  DFF_X1 \DRAM_mem_reg[10][2]  ( .D(n8917), .CK(CLK), .Q(n6476), .QN(n37616)
         );
  DFF_X1 \DRAM_mem_reg[10][1]  ( .D(n8916), .CK(CLK), .Q(n6475), .QN(n37615)
         );
  DFF_X1 \DRAM_mem_reg[10][0]  ( .D(n8915), .CK(CLK), .Q(n6474), .QN(n37614)
         );
  DFF_X1 \DRAM_mem_reg[11][31]  ( .D(n8914), .CK(CLK), .Q(n5560), .QN(n37485)
         );
  DFF_X1 \DRAM_mem_reg[11][30]  ( .D(n8913), .CK(CLK), .Q(n5610), .QN(n37484)
         );
  DFF_X1 \DRAM_mem_reg[11][29]  ( .D(n8912), .CK(CLK), .Q(n5652), .QN(n37483)
         );
  DFF_X1 \DRAM_mem_reg[11][28]  ( .D(n8911), .CK(CLK), .Q(n5694), .QN(n37482)
         );
  DFF_X1 \DRAM_mem_reg[11][27]  ( .D(n8910), .CK(CLK), .Q(n5736), .QN(n37481)
         );
  DFF_X1 \DRAM_mem_reg[11][26]  ( .D(n8909), .CK(CLK), .Q(n5778), .QN(n37480)
         );
  DFF_X1 \DRAM_mem_reg[11][25]  ( .D(n8908), .CK(CLK), .Q(n5820), .QN(n37479)
         );
  DFF_X1 \DRAM_mem_reg[11][24]  ( .D(n8907), .CK(CLK), .Q(n5862), .QN(n37478)
         );
  DFF_X1 \DRAM_mem_reg[11][23]  ( .D(n8906), .CK(CLK), .Q(n5904), .QN(n37477)
         );
  DFF_X1 \DRAM_mem_reg[11][22]  ( .D(n8905), .CK(CLK), .Q(n5946), .QN(n37476)
         );
  DFF_X1 \DRAM_mem_reg[11][21]  ( .D(n8904), .CK(CLK), .Q(n5988), .QN(n37475)
         );
  DFF_X1 \DRAM_mem_reg[11][20]  ( .D(n8903), .CK(CLK), .Q(n6030), .QN(n37474)
         );
  DFF_X1 \DRAM_mem_reg[11][19]  ( .D(n8902), .CK(CLK), .Q(n6072), .QN(n37473)
         );
  DFF_X1 \DRAM_mem_reg[11][18]  ( .D(n8901), .CK(CLK), .Q(n6114), .QN(n37472)
         );
  DFF_X1 \DRAM_mem_reg[11][17]  ( .D(n8900), .CK(CLK), .Q(n6156), .QN(n37471)
         );
  DFF_X1 \DRAM_mem_reg[11][16]  ( .D(n8899), .CK(CLK), .Q(n6198), .QN(n37470)
         );
  DFF_X1 \DRAM_mem_reg[11][15]  ( .D(n8898), .CK(CLK), .Q(n6240), .QN(n37469)
         );
  DFF_X1 \DRAM_mem_reg[11][14]  ( .D(n8897), .CK(CLK), .Q(n6282), .QN(n37468)
         );
  DFF_X1 \DRAM_mem_reg[11][13]  ( .D(n8896), .CK(CLK), .Q(n6324), .QN(n37467)
         );
  DFF_X1 \DRAM_mem_reg[11][12]  ( .D(n8895), .CK(CLK), .Q(n6366), .QN(n37466)
         );
  DFF_X1 \DRAM_mem_reg[11][11]  ( .D(n8894), .CK(CLK), .Q(n6536), .QN(n37465)
         );
  DFF_X1 \DRAM_mem_reg[11][10]  ( .D(n8893), .CK(CLK), .Q(n6578), .QN(n37464)
         );
  DFF_X1 \DRAM_mem_reg[11][9]  ( .D(n8892), .CK(CLK), .Q(n6620), .QN(n37463)
         );
  DFF_X1 \DRAM_mem_reg[11][8]  ( .D(n8891), .CK(CLK), .Q(n6662), .QN(n37462)
         );
  DFF_X1 \DRAM_mem_reg[11][7]  ( .D(n8890), .CK(CLK), .Q(n9296), .QN(n37461)
         );
  DFF_X1 \DRAM_mem_reg[11][6]  ( .D(n8889), .CK(CLK), .Q(n9338), .QN(n37460)
         );
  DFF_X1 \DRAM_mem_reg[11][5]  ( .D(n8888), .CK(CLK), .Q(n9380), .QN(n37459)
         );
  DFF_X1 \DRAM_mem_reg[11][4]  ( .D(n8887), .CK(CLK), .Q(n9422), .QN(n37458)
         );
  DFF_X1 \DRAM_mem_reg[11][3]  ( .D(n8886), .CK(CLK), .Q(n9464), .QN(n37457)
         );
  DFF_X1 \DRAM_mem_reg[11][2]  ( .D(n8885), .CK(CLK), .Q(n9506), .QN(n37456)
         );
  DFF_X1 \DRAM_mem_reg[11][1]  ( .D(n8884), .CK(CLK), .Q(n9548), .QN(n37455)
         );
  DFF_X1 \DRAM_mem_reg[11][0]  ( .D(n8883), .CK(CLK), .Q(n9613), .QN(n37454)
         );
  DFF_X1 \DRAM_mem_reg[12][31]  ( .D(n8882), .CK(CLK), .QN(n35701) );
  DFF_X1 \DRAM_mem_reg[12][30]  ( .D(n8881), .CK(CLK), .QN(n35700) );
  DFF_X1 \DRAM_mem_reg[12][29]  ( .D(n8880), .CK(CLK), .QN(n35699) );
  DFF_X1 \DRAM_mem_reg[12][28]  ( .D(n8879), .CK(CLK), .QN(n35698) );
  DFF_X1 \DRAM_mem_reg[12][27]  ( .D(n8878), .CK(CLK), .QN(n35697) );
  DFF_X1 \DRAM_mem_reg[12][26]  ( .D(n8877), .CK(CLK), .QN(n35696) );
  DFF_X1 \DRAM_mem_reg[12][25]  ( .D(n8876), .CK(CLK), .QN(n35695) );
  DFF_X1 \DRAM_mem_reg[12][24]  ( .D(n8875), .CK(CLK), .QN(n35694) );
  DFF_X1 \DRAM_mem_reg[12][23]  ( .D(n8874), .CK(CLK), .QN(n35829) );
  DFF_X1 \DRAM_mem_reg[12][22]  ( .D(n8873), .CK(CLK), .QN(n35828) );
  DFF_X1 \DRAM_mem_reg[12][21]  ( .D(n8872), .CK(CLK), .QN(n35827) );
  DFF_X1 \DRAM_mem_reg[12][20]  ( .D(n8871), .CK(CLK), .QN(n35826) );
  DFF_X1 \DRAM_mem_reg[12][19]  ( .D(n8870), .CK(CLK), .QN(n35825) );
  DFF_X1 \DRAM_mem_reg[12][18]  ( .D(n8869), .CK(CLK), .QN(n35824) );
  DFF_X1 \DRAM_mem_reg[12][17]  ( .D(n8868), .CK(CLK), .QN(n35823) );
  DFF_X1 \DRAM_mem_reg[12][16]  ( .D(n8867), .CK(CLK), .QN(n35822) );
  DFF_X1 \DRAM_mem_reg[12][15]  ( .D(n8866), .CK(CLK), .QN(n35821) );
  DFF_X1 \DRAM_mem_reg[12][14]  ( .D(n8865), .CK(CLK), .QN(n35820) );
  DFF_X1 \DRAM_mem_reg[12][13]  ( .D(n8864), .CK(CLK), .QN(n35819) );
  DFF_X1 \DRAM_mem_reg[12][12]  ( .D(n8863), .CK(CLK), .QN(n35818) );
  DFF_X1 \DRAM_mem_reg[12][11]  ( .D(n8862), .CK(CLK), .QN(n35817) );
  DFF_X1 \DRAM_mem_reg[12][10]  ( .D(n8861), .CK(CLK), .QN(n35816) );
  DFF_X1 \DRAM_mem_reg[12][9]  ( .D(n8860), .CK(CLK), .QN(n35815) );
  DFF_X1 \DRAM_mem_reg[12][8]  ( .D(n8859), .CK(CLK), .QN(n35814) );
  DFF_X1 \DRAM_mem_reg[12][7]  ( .D(n8858), .CK(CLK), .QN(n35813) );
  DFF_X1 \DRAM_mem_reg[12][6]  ( .D(n8857), .CK(CLK), .QN(n35812) );
  DFF_X1 \DRAM_mem_reg[12][5]  ( .D(n8856), .CK(CLK), .QN(n35811) );
  DFF_X1 \DRAM_mem_reg[12][4]  ( .D(n8855), .CK(CLK), .QN(n35810) );
  DFF_X1 \DRAM_mem_reg[12][3]  ( .D(n8854), .CK(CLK), .QN(n35809) );
  DFF_X1 \DRAM_mem_reg[12][2]  ( .D(n8853), .CK(CLK), .QN(n35808) );
  DFF_X1 \DRAM_mem_reg[12][1]  ( .D(n8852), .CK(CLK), .QN(n35807) );
  DFF_X1 \DRAM_mem_reg[12][0]  ( .D(n8851), .CK(CLK), .QN(n35806) );
  DFF_X1 \DRAM_mem_reg[13][31]  ( .D(n8850), .CK(CLK), .QN(n36213) );
  DFF_X1 \DRAM_mem_reg[13][30]  ( .D(n8849), .CK(CLK), .QN(n36212) );
  DFF_X1 \DRAM_mem_reg[13][29]  ( .D(n8848), .CK(CLK), .QN(n36211) );
  DFF_X1 \DRAM_mem_reg[13][28]  ( .D(n8847), .CK(CLK), .QN(n36210) );
  DFF_X1 \DRAM_mem_reg[13][27]  ( .D(n8846), .CK(CLK), .QN(n36209) );
  DFF_X1 \DRAM_mem_reg[13][26]  ( .D(n8845), .CK(CLK), .QN(n36208) );
  DFF_X1 \DRAM_mem_reg[13][25]  ( .D(n8844), .CK(CLK), .QN(n36207) );
  DFF_X1 \DRAM_mem_reg[13][24]  ( .D(n8843), .CK(CLK), .QN(n36206) );
  DFF_X1 \DRAM_mem_reg[13][23]  ( .D(n8842), .CK(CLK), .QN(n36341) );
  DFF_X1 \DRAM_mem_reg[13][22]  ( .D(n8841), .CK(CLK), .QN(n36340) );
  DFF_X1 \DRAM_mem_reg[13][21]  ( .D(n8840), .CK(CLK), .QN(n36339) );
  DFF_X1 \DRAM_mem_reg[13][20]  ( .D(n8839), .CK(CLK), .QN(n36338) );
  DFF_X1 \DRAM_mem_reg[13][19]  ( .D(n8838), .CK(CLK), .QN(n36337) );
  DFF_X1 \DRAM_mem_reg[13][18]  ( .D(n8837), .CK(CLK), .QN(n36336) );
  DFF_X1 \DRAM_mem_reg[13][17]  ( .D(n8836), .CK(CLK), .QN(n36335) );
  DFF_X1 \DRAM_mem_reg[13][16]  ( .D(n8835), .CK(CLK), .QN(n36334) );
  DFF_X1 \DRAM_mem_reg[13][15]  ( .D(n8834), .CK(CLK), .QN(n36333) );
  DFF_X1 \DRAM_mem_reg[13][14]  ( .D(n8833), .CK(CLK), .QN(n36332) );
  DFF_X1 \DRAM_mem_reg[13][13]  ( .D(n8832), .CK(CLK), .QN(n36331) );
  DFF_X1 \DRAM_mem_reg[13][12]  ( .D(n8831), .CK(CLK), .QN(n36330) );
  DFF_X1 \DRAM_mem_reg[13][11]  ( .D(n8830), .CK(CLK), .QN(n36329) );
  DFF_X1 \DRAM_mem_reg[13][10]  ( .D(n8829), .CK(CLK), .QN(n36328) );
  DFF_X1 \DRAM_mem_reg[13][9]  ( .D(n8828), .CK(CLK), .QN(n36327) );
  DFF_X1 \DRAM_mem_reg[13][8]  ( .D(n8827), .CK(CLK), .QN(n36326) );
  DFF_X1 \DRAM_mem_reg[13][7]  ( .D(n8826), .CK(CLK), .QN(n36325) );
  DFF_X1 \DRAM_mem_reg[13][6]  ( .D(n8825), .CK(CLK), .QN(n36324) );
  DFF_X1 \DRAM_mem_reg[13][5]  ( .D(n8824), .CK(CLK), .QN(n36323) );
  DFF_X1 \DRAM_mem_reg[13][4]  ( .D(n8823), .CK(CLK), .QN(n36322) );
  DFF_X1 \DRAM_mem_reg[13][3]  ( .D(n8822), .CK(CLK), .QN(n36321) );
  DFF_X1 \DRAM_mem_reg[13][2]  ( .D(n8821), .CK(CLK), .QN(n36320) );
  DFF_X1 \DRAM_mem_reg[13][1]  ( .D(n8820), .CK(CLK), .QN(n36319) );
  DFF_X1 \DRAM_mem_reg[13][0]  ( .D(n8819), .CK(CLK), .QN(n36318) );
  DFF_X1 \DRAM_mem_reg[14][31]  ( .D(n8818), .CK(CLK), .QN(n35189) );
  DFF_X1 \DRAM_mem_reg[14][30]  ( .D(n8817), .CK(CLK), .QN(n35188) );
  DFF_X1 \DRAM_mem_reg[14][29]  ( .D(n8816), .CK(CLK), .QN(n35187) );
  DFF_X1 \DRAM_mem_reg[14][28]  ( .D(n8815), .CK(CLK), .QN(n35186) );
  DFF_X1 \DRAM_mem_reg[14][27]  ( .D(n8814), .CK(CLK), .QN(n35185) );
  DFF_X1 \DRAM_mem_reg[14][26]  ( .D(n8813), .CK(CLK), .QN(n35184) );
  DFF_X1 \DRAM_mem_reg[14][25]  ( .D(n8812), .CK(CLK), .QN(n35183) );
  DFF_X1 \DRAM_mem_reg[14][24]  ( .D(n8811), .CK(CLK), .QN(n35182) );
  DFF_X1 \DRAM_mem_reg[14][23]  ( .D(n8810), .CK(CLK), .QN(n35317) );
  DFF_X1 \DRAM_mem_reg[14][22]  ( .D(n8809), .CK(CLK), .QN(n35316) );
  DFF_X1 \DRAM_mem_reg[14][21]  ( .D(n8808), .CK(CLK), .QN(n35315) );
  DFF_X1 \DRAM_mem_reg[14][20]  ( .D(n8807), .CK(CLK), .QN(n35314) );
  DFF_X1 \DRAM_mem_reg[14][19]  ( .D(n8806), .CK(CLK), .QN(n35313) );
  DFF_X1 \DRAM_mem_reg[14][18]  ( .D(n8805), .CK(CLK), .QN(n35312) );
  DFF_X1 \DRAM_mem_reg[14][17]  ( .D(n8804), .CK(CLK), .QN(n35311) );
  DFF_X1 \DRAM_mem_reg[14][16]  ( .D(n8803), .CK(CLK), .QN(n35310) );
  DFF_X1 \DRAM_mem_reg[14][15]  ( .D(n8802), .CK(CLK), .QN(n35309) );
  DFF_X1 \DRAM_mem_reg[14][14]  ( .D(n8801), .CK(CLK), .QN(n35308) );
  DFF_X1 \DRAM_mem_reg[14][13]  ( .D(n8800), .CK(CLK), .QN(n35307) );
  DFF_X1 \DRAM_mem_reg[14][12]  ( .D(n8799), .CK(CLK), .QN(n35306) );
  DFF_X1 \DRAM_mem_reg[14][11]  ( .D(n8798), .CK(CLK), .QN(n35305) );
  DFF_X1 \DRAM_mem_reg[14][10]  ( .D(n8797), .CK(CLK), .QN(n35304) );
  DFF_X1 \DRAM_mem_reg[14][9]  ( .D(n8796), .CK(CLK), .QN(n35303) );
  DFF_X1 \DRAM_mem_reg[14][8]  ( .D(n8795), .CK(CLK), .QN(n35302) );
  DFF_X1 \DRAM_mem_reg[14][7]  ( .D(n8794), .CK(CLK), .QN(n35301) );
  DFF_X1 \DRAM_mem_reg[14][6]  ( .D(n8793), .CK(CLK), .QN(n35300) );
  DFF_X1 \DRAM_mem_reg[14][5]  ( .D(n8792), .CK(CLK), .QN(n35299) );
  DFF_X1 \DRAM_mem_reg[14][4]  ( .D(n8791), .CK(CLK), .QN(n35298) );
  DFF_X1 \DRAM_mem_reg[14][3]  ( .D(n8790), .CK(CLK), .QN(n35297) );
  DFF_X1 \DRAM_mem_reg[14][2]  ( .D(n8789), .CK(CLK), .QN(n35296) );
  DFF_X1 \DRAM_mem_reg[14][1]  ( .D(n8788), .CK(CLK), .QN(n35295) );
  DFF_X1 \DRAM_mem_reg[14][0]  ( .D(n8787), .CK(CLK), .QN(n35294) );
  DFF_X1 \DRAM_mem_reg[15][31]  ( .D(n8786), .CK(CLK), .Q(n6473), .QN(n37613)
         );
  DFF_X1 \DRAM_mem_reg[15][30]  ( .D(n8785), .CK(CLK), .Q(n6472), .QN(n37612)
         );
  DFF_X1 \DRAM_mem_reg[15][29]  ( .D(n8784), .CK(CLK), .Q(n6471), .QN(n37611)
         );
  DFF_X1 \DRAM_mem_reg[15][28]  ( .D(n8783), .CK(CLK), .Q(n6470), .QN(n37610)
         );
  DFF_X1 \DRAM_mem_reg[15][27]  ( .D(n8782), .CK(CLK), .Q(n6469), .QN(n37609)
         );
  DFF_X1 \DRAM_mem_reg[15][26]  ( .D(n8781), .CK(CLK), .Q(n6468), .QN(n37608)
         );
  DFF_X1 \DRAM_mem_reg[15][25]  ( .D(n8780), .CK(CLK), .Q(n6467), .QN(n37607)
         );
  DFF_X1 \DRAM_mem_reg[15][24]  ( .D(n8779), .CK(CLK), .Q(n6466), .QN(n37606)
         );
  DFF_X1 \DRAM_mem_reg[15][23]  ( .D(n8778), .CK(CLK), .Q(n6465), .QN(n37605)
         );
  DFF_X1 \DRAM_mem_reg[15][22]  ( .D(n8777), .CK(CLK), .Q(n6464), .QN(n37604)
         );
  DFF_X1 \DRAM_mem_reg[15][21]  ( .D(n8776), .CK(CLK), .Q(n6463), .QN(n37603)
         );
  DFF_X1 \DRAM_mem_reg[15][20]  ( .D(n8775), .CK(CLK), .Q(n6462), .QN(n37602)
         );
  DFF_X1 \DRAM_mem_reg[15][19]  ( .D(n8774), .CK(CLK), .Q(n6461), .QN(n37601)
         );
  DFF_X1 \DRAM_mem_reg[15][18]  ( .D(n8773), .CK(CLK), .Q(n6460), .QN(n37600)
         );
  DFF_X1 \DRAM_mem_reg[15][17]  ( .D(n8772), .CK(CLK), .Q(n6459), .QN(n37599)
         );
  DFF_X1 \DRAM_mem_reg[15][16]  ( .D(n8771), .CK(CLK), .Q(n6458), .QN(n37598)
         );
  DFF_X1 \DRAM_mem_reg[15][15]  ( .D(n8770), .CK(CLK), .Q(n6457), .QN(n37597)
         );
  DFF_X1 \DRAM_mem_reg[15][14]  ( .D(n8769), .CK(CLK), .Q(n6456), .QN(n37596)
         );
  DFF_X1 \DRAM_mem_reg[15][13]  ( .D(n8768), .CK(CLK), .Q(n6455), .QN(n37595)
         );
  DFF_X1 \DRAM_mem_reg[15][12]  ( .D(n8767), .CK(CLK), .Q(n6454), .QN(n37594)
         );
  DFF_X1 \DRAM_mem_reg[15][11]  ( .D(n8766), .CK(CLK), .Q(n6453), .QN(n37593)
         );
  DFF_X1 \DRAM_mem_reg[15][10]  ( .D(n8765), .CK(CLK), .Q(n6452), .QN(n37592)
         );
  DFF_X1 \DRAM_mem_reg[15][9]  ( .D(n8764), .CK(CLK), .Q(n6451), .QN(n37591)
         );
  DFF_X1 \DRAM_mem_reg[15][8]  ( .D(n8763), .CK(CLK), .Q(n6450), .QN(n37590)
         );
  DFF_X1 \DRAM_mem_reg[15][7]  ( .D(n8762), .CK(CLK), .Q(n6448), .QN(n37589)
         );
  DFF_X1 \DRAM_mem_reg[15][6]  ( .D(n8761), .CK(CLK), .Q(n6445), .QN(n37588)
         );
  DFF_X1 \DRAM_mem_reg[15][5]  ( .D(n8760), .CK(CLK), .Q(n6442), .QN(n37587)
         );
  DFF_X1 \DRAM_mem_reg[15][4]  ( .D(n8759), .CK(CLK), .Q(n6440), .QN(n37586)
         );
  DFF_X1 \DRAM_mem_reg[15][3]  ( .D(n8758), .CK(CLK), .Q(n6439), .QN(n37585)
         );
  DFF_X1 \DRAM_mem_reg[15][2]  ( .D(n8757), .CK(CLK), .Q(n6438), .QN(n37584)
         );
  DFF_X1 \DRAM_mem_reg[15][1]  ( .D(n8756), .CK(CLK), .Q(n6437), .QN(n37583)
         );
  DFF_X1 \DRAM_mem_reg[15][0]  ( .D(n8755), .CK(CLK), .Q(n6436), .QN(n37582)
         );
  DFF_X1 \DRAM_mem_reg[16][31]  ( .D(n8754), .CK(CLK), .QN(n35181) );
  DFF_X1 \DRAM_mem_reg[16][30]  ( .D(n8753), .CK(CLK), .QN(n35180) );
  DFF_X1 \DRAM_mem_reg[16][29]  ( .D(n8752), .CK(CLK), .QN(n35179) );
  DFF_X1 \DRAM_mem_reg[16][28]  ( .D(n8751), .CK(CLK), .QN(n35178) );
  DFF_X1 \DRAM_mem_reg[16][27]  ( .D(n8750), .CK(CLK), .QN(n35177) );
  DFF_X1 \DRAM_mem_reg[16][26]  ( .D(n8749), .CK(CLK), .QN(n35176) );
  DFF_X1 \DRAM_mem_reg[16][25]  ( .D(n8748), .CK(CLK), .QN(n35175) );
  DFF_X1 \DRAM_mem_reg[16][24]  ( .D(n8747), .CK(CLK), .QN(n35174) );
  DFF_X1 \DRAM_mem_reg[16][23]  ( .D(n8746), .CK(CLK), .QN(n35293) );
  DFF_X1 \DRAM_mem_reg[16][22]  ( .D(n8745), .CK(CLK), .QN(n35292) );
  DFF_X1 \DRAM_mem_reg[16][21]  ( .D(n8744), .CK(CLK), .QN(n35291) );
  DFF_X1 \DRAM_mem_reg[16][20]  ( .D(n8743), .CK(CLK), .QN(n35290) );
  DFF_X1 \DRAM_mem_reg[16][19]  ( .D(n8742), .CK(CLK), .QN(n35289) );
  DFF_X1 \DRAM_mem_reg[16][18]  ( .D(n8741), .CK(CLK), .QN(n35288) );
  DFF_X1 \DRAM_mem_reg[16][17]  ( .D(n8740), .CK(CLK), .QN(n35287) );
  DFF_X1 \DRAM_mem_reg[16][16]  ( .D(n8739), .CK(CLK), .QN(n35286) );
  DFF_X1 \DRAM_mem_reg[16][15]  ( .D(n8738), .CK(CLK), .QN(n35285) );
  DFF_X1 \DRAM_mem_reg[16][14]  ( .D(n8737), .CK(CLK), .QN(n35284) );
  DFF_X1 \DRAM_mem_reg[16][13]  ( .D(n8736), .CK(CLK), .QN(n35283) );
  DFF_X1 \DRAM_mem_reg[16][12]  ( .D(n8735), .CK(CLK), .QN(n35282) );
  DFF_X1 \DRAM_mem_reg[16][11]  ( .D(n8734), .CK(CLK), .QN(n35281) );
  DFF_X1 \DRAM_mem_reg[16][10]  ( .D(n8733), .CK(CLK), .QN(n35280) );
  DFF_X1 \DRAM_mem_reg[16][9]  ( .D(n8732), .CK(CLK), .QN(n35279) );
  DFF_X1 \DRAM_mem_reg[16][8]  ( .D(n8731), .CK(CLK), .QN(n35278) );
  DFF_X1 \DRAM_mem_reg[16][7]  ( .D(n8730), .CK(CLK), .QN(n35277) );
  DFF_X1 \DRAM_mem_reg[16][6]  ( .D(n8729), .CK(CLK), .QN(n35276) );
  DFF_X1 \DRAM_mem_reg[16][5]  ( .D(n8728), .CK(CLK), .QN(n35275) );
  DFF_X1 \DRAM_mem_reg[16][4]  ( .D(n8727), .CK(CLK), .QN(n35274) );
  DFF_X1 \DRAM_mem_reg[16][3]  ( .D(n8726), .CK(CLK), .QN(n35273) );
  DFF_X1 \DRAM_mem_reg[16][2]  ( .D(n8725), .CK(CLK), .QN(n35272) );
  DFF_X1 \DRAM_mem_reg[16][1]  ( .D(n8724), .CK(CLK), .QN(n35271) );
  DFF_X1 \DRAM_mem_reg[16][0]  ( .D(n8723), .CK(CLK), .QN(n35270) );
  DFF_X1 \DRAM_mem_reg[17][31]  ( .D(n8722), .CK(CLK), .QN(n35693) );
  DFF_X1 \DRAM_mem_reg[17][30]  ( .D(n8721), .CK(CLK), .QN(n35692) );
  DFF_X1 \DRAM_mem_reg[17][29]  ( .D(n8720), .CK(CLK), .QN(n35691) );
  DFF_X1 \DRAM_mem_reg[17][28]  ( .D(n8719), .CK(CLK), .QN(n35690) );
  DFF_X1 \DRAM_mem_reg[17][27]  ( .D(n8718), .CK(CLK), .QN(n35689) );
  DFF_X1 \DRAM_mem_reg[17][26]  ( .D(n8717), .CK(CLK), .QN(n35688) );
  DFF_X1 \DRAM_mem_reg[17][25]  ( .D(n8716), .CK(CLK), .QN(n35687) );
  DFF_X1 \DRAM_mem_reg[17][24]  ( .D(n8715), .CK(CLK), .QN(n35686) );
  DFF_X1 \DRAM_mem_reg[17][23]  ( .D(n8714), .CK(CLK), .QN(n35805) );
  DFF_X1 \DRAM_mem_reg[17][22]  ( .D(n8713), .CK(CLK), .QN(n35804) );
  DFF_X1 \DRAM_mem_reg[17][21]  ( .D(n8712), .CK(CLK), .QN(n35803) );
  DFF_X1 \DRAM_mem_reg[17][20]  ( .D(n8711), .CK(CLK), .QN(n35802) );
  DFF_X1 \DRAM_mem_reg[17][19]  ( .D(n8710), .CK(CLK), .QN(n35801) );
  DFF_X1 \DRAM_mem_reg[17][18]  ( .D(n8709), .CK(CLK), .QN(n35800) );
  DFF_X1 \DRAM_mem_reg[17][17]  ( .D(n8708), .CK(CLK), .QN(n35799) );
  DFF_X1 \DRAM_mem_reg[17][16]  ( .D(n8707), .CK(CLK), .QN(n35798) );
  DFF_X1 \DRAM_mem_reg[17][15]  ( .D(n8706), .CK(CLK), .QN(n35797) );
  DFF_X1 \DRAM_mem_reg[17][14]  ( .D(n8705), .CK(CLK), .QN(n35796) );
  DFF_X1 \DRAM_mem_reg[17][13]  ( .D(n8704), .CK(CLK), .QN(n35795) );
  DFF_X1 \DRAM_mem_reg[17][12]  ( .D(n8703), .CK(CLK), .QN(n35794) );
  DFF_X1 \DRAM_mem_reg[17][11]  ( .D(n8702), .CK(CLK), .QN(n35793) );
  DFF_X1 \DRAM_mem_reg[17][10]  ( .D(n8701), .CK(CLK), .QN(n35792) );
  DFF_X1 \DRAM_mem_reg[17][9]  ( .D(n8700), .CK(CLK), .QN(n35791) );
  DFF_X1 \DRAM_mem_reg[17][8]  ( .D(n8699), .CK(CLK), .QN(n35790) );
  DFF_X1 \DRAM_mem_reg[17][7]  ( .D(n8698), .CK(CLK), .QN(n35789) );
  DFF_X1 \DRAM_mem_reg[17][6]  ( .D(n8697), .CK(CLK), .QN(n35788) );
  DFF_X1 \DRAM_mem_reg[17][5]  ( .D(n8696), .CK(CLK), .QN(n35787) );
  DFF_X1 \DRAM_mem_reg[17][4]  ( .D(n8695), .CK(CLK), .QN(n35786) );
  DFF_X1 \DRAM_mem_reg[17][3]  ( .D(n8694), .CK(CLK), .QN(n35785) );
  DFF_X1 \DRAM_mem_reg[17][2]  ( .D(n8693), .CK(CLK), .QN(n35784) );
  DFF_X1 \DRAM_mem_reg[17][1]  ( .D(n8692), .CK(CLK), .QN(n35783) );
  DFF_X1 \DRAM_mem_reg[17][0]  ( .D(n8691), .CK(CLK), .QN(n35782) );
  DFF_X1 \DRAM_mem_reg[18][31]  ( .D(n8690), .CK(CLK), .Q(net254318), .QN(
        n37165) );
  DFF_X1 \DRAM_mem_reg[18][30]  ( .D(n8689), .CK(CLK), .Q(net254317), .QN(
        n37164) );
  DFF_X1 \DRAM_mem_reg[18][29]  ( .D(n8688), .CK(CLK), .Q(net254316), .QN(
        n37163) );
  DFF_X1 \DRAM_mem_reg[18][28]  ( .D(n8687), .CK(CLK), .Q(net254315), .QN(
        n37162) );
  DFF_X1 \DRAM_mem_reg[18][27]  ( .D(n8686), .CK(CLK), .Q(net254314), .QN(
        n37161) );
  DFF_X1 \DRAM_mem_reg[18][26]  ( .D(n8685), .CK(CLK), .Q(net254313), .QN(
        n37160) );
  DFF_X1 \DRAM_mem_reg[18][25]  ( .D(n8684), .CK(CLK), .Q(net254312), .QN(
        n37159) );
  DFF_X1 \DRAM_mem_reg[18][24]  ( .D(n8683), .CK(CLK), .Q(net254311), .QN(
        n37158) );
  DFF_X1 \DRAM_mem_reg[18][23]  ( .D(n8682), .CK(CLK), .Q(net254310), .QN(
        n37453) );
  DFF_X1 \DRAM_mem_reg[18][22]  ( .D(n8681), .CK(CLK), .Q(net254309), .QN(
        n37452) );
  DFF_X1 \DRAM_mem_reg[18][21]  ( .D(n8680), .CK(CLK), .Q(net254308), .QN(
        n37451) );
  DFF_X1 \DRAM_mem_reg[18][20]  ( .D(n8679), .CK(CLK), .Q(net254307), .QN(
        n37450) );
  DFF_X1 \DRAM_mem_reg[18][19]  ( .D(n8678), .CK(CLK), .Q(net254306), .QN(
        n37449) );
  DFF_X1 \DRAM_mem_reg[18][18]  ( .D(n8677), .CK(CLK), .Q(net254305), .QN(
        n37448) );
  DFF_X1 \DRAM_mem_reg[18][17]  ( .D(n8676), .CK(CLK), .Q(net254304), .QN(
        n37447) );
  DFF_X1 \DRAM_mem_reg[18][16]  ( .D(n8675), .CK(CLK), .Q(net254303), .QN(
        n37446) );
  DFF_X1 \DRAM_mem_reg[18][15]  ( .D(n8674), .CK(CLK), .Q(net254302), .QN(
        n37445) );
  DFF_X1 \DRAM_mem_reg[18][14]  ( .D(n8673), .CK(CLK), .Q(net254301), .QN(
        n37444) );
  DFF_X1 \DRAM_mem_reg[18][13]  ( .D(n8672), .CK(CLK), .Q(net254300), .QN(
        n37443) );
  DFF_X1 \DRAM_mem_reg[18][12]  ( .D(n8671), .CK(CLK), .Q(net254299), .QN(
        n37442) );
  DFF_X1 \DRAM_mem_reg[18][11]  ( .D(n8670), .CK(CLK), .Q(net254298), .QN(
        n37441) );
  DFF_X1 \DRAM_mem_reg[18][10]  ( .D(n8669), .CK(CLK), .Q(net254297), .QN(
        n37440) );
  DFF_X1 \DRAM_mem_reg[18][9]  ( .D(n8668), .CK(CLK), .Q(net254296), .QN(
        n37439) );
  DFF_X1 \DRAM_mem_reg[18][8]  ( .D(n8667), .CK(CLK), .Q(net254295), .QN(
        n37438) );
  DFF_X1 \DRAM_mem_reg[18][7]  ( .D(n8666), .CK(CLK), .Q(net254294), .QN(
        n37437) );
  DFF_X1 \DRAM_mem_reg[18][6]  ( .D(n8665), .CK(CLK), .Q(net254293), .QN(
        n37436) );
  DFF_X1 \DRAM_mem_reg[18][5]  ( .D(n8664), .CK(CLK), .Q(net254292), .QN(
        n37435) );
  DFF_X1 \DRAM_mem_reg[18][4]  ( .D(n8663), .CK(CLK), .Q(net254291), .QN(
        n37434) );
  DFF_X1 \DRAM_mem_reg[18][3]  ( .D(n8662), .CK(CLK), .Q(net254290), .QN(
        n37433) );
  DFF_X1 \DRAM_mem_reg[18][2]  ( .D(n8661), .CK(CLK), .Q(net254289), .QN(
        n37432) );
  DFF_X1 \DRAM_mem_reg[18][1]  ( .D(n8660), .CK(CLK), .Q(net254288), .QN(
        n37431) );
  DFF_X1 \DRAM_mem_reg[18][0]  ( .D(n8659), .CK(CLK), .Q(net254287), .QN(
        n37430) );
  DFF_X1 \DRAM_mem_reg[19][31]  ( .D(n8658), .CK(CLK), .QN(n36435) );
  DFF_X1 \DRAM_mem_reg[19][30]  ( .D(n8657), .CK(CLK), .QN(n36426) );
  DFF_X1 \DRAM_mem_reg[19][29]  ( .D(n8656), .CK(CLK), .QN(n36417) );
  DFF_X1 \DRAM_mem_reg[19][28]  ( .D(n8655), .CK(CLK), .QN(n36408) );
  DFF_X1 \DRAM_mem_reg[19][27]  ( .D(n8654), .CK(CLK), .QN(n36399) );
  DFF_X1 \DRAM_mem_reg[19][26]  ( .D(n8653), .CK(CLK), .QN(n36390) );
  DFF_X1 \DRAM_mem_reg[19][25]  ( .D(n8652), .CK(CLK), .QN(n36381) );
  DFF_X1 \DRAM_mem_reg[19][24]  ( .D(n8651), .CK(CLK), .QN(n36372) );
  DFF_X1 \DRAM_mem_reg[19][23]  ( .D(n8650), .CK(CLK), .QN(n36589) );
  DFF_X1 \DRAM_mem_reg[19][22]  ( .D(n8649), .CK(CLK), .QN(n36587) );
  DFF_X1 \DRAM_mem_reg[19][21]  ( .D(n8648), .CK(CLK), .QN(n36585) );
  DFF_X1 \DRAM_mem_reg[19][20]  ( .D(n8647), .CK(CLK), .QN(n36583) );
  DFF_X1 \DRAM_mem_reg[19][19]  ( .D(n8646), .CK(CLK), .QN(n36581) );
  DFF_X1 \DRAM_mem_reg[19][18]  ( .D(n8645), .CK(CLK), .QN(n36579) );
  DFF_X1 \DRAM_mem_reg[19][17]  ( .D(n8644), .CK(CLK), .QN(n36577) );
  DFF_X1 \DRAM_mem_reg[19][16]  ( .D(n8643), .CK(CLK), .QN(n36575) );
  DFF_X1 \DRAM_mem_reg[19][15]  ( .D(n8642), .CK(CLK), .QN(n36573) );
  DFF_X1 \DRAM_mem_reg[19][14]  ( .D(n8641), .CK(CLK), .QN(n36571) );
  DFF_X1 \DRAM_mem_reg[19][13]  ( .D(n8640), .CK(CLK), .QN(n36569) );
  DFF_X1 \DRAM_mem_reg[19][12]  ( .D(n8639), .CK(CLK), .QN(n36567) );
  DFF_X1 \DRAM_mem_reg[19][11]  ( .D(n8638), .CK(CLK), .QN(n36565) );
  DFF_X1 \DRAM_mem_reg[19][10]  ( .D(n8637), .CK(CLK), .QN(n36563) );
  DFF_X1 \DRAM_mem_reg[19][9]  ( .D(n8636), .CK(CLK), .QN(n36561) );
  DFF_X1 \DRAM_mem_reg[19][8]  ( .D(n8635), .CK(CLK), .QN(n36559) );
  DFF_X1 \DRAM_mem_reg[19][7]  ( .D(n8634), .CK(CLK), .QN(n36557) );
  DFF_X1 \DRAM_mem_reg[19][6]  ( .D(n8633), .CK(CLK), .QN(n36555) );
  DFF_X1 \DRAM_mem_reg[19][5]  ( .D(n8632), .CK(CLK), .QN(n36553) );
  DFF_X1 \DRAM_mem_reg[19][4]  ( .D(n8631), .CK(CLK), .QN(n36551) );
  DFF_X1 \DRAM_mem_reg[19][3]  ( .D(n8630), .CK(CLK), .QN(n36549) );
  DFF_X1 \DRAM_mem_reg[19][2]  ( .D(n8629), .CK(CLK), .QN(n36547) );
  DFF_X1 \DRAM_mem_reg[19][1]  ( .D(n8628), .CK(CLK), .QN(n36545) );
  DFF_X1 \DRAM_mem_reg[19][0]  ( .D(n8627), .CK(CLK), .QN(n36543) );
  DFF_X1 \DRAM_mem_reg[20][31]  ( .D(n8626), .CK(CLK), .Q(net254286), .QN(
        n36781) );
  DFF_X1 \DRAM_mem_reg[20][30]  ( .D(n8625), .CK(CLK), .Q(net254285), .QN(
        n36780) );
  DFF_X1 \DRAM_mem_reg[20][29]  ( .D(n8624), .CK(CLK), .Q(net254284), .QN(
        n36779) );
  DFF_X1 \DRAM_mem_reg[20][28]  ( .D(n8623), .CK(CLK), .Q(net254283), .QN(
        n36778) );
  DFF_X1 \DRAM_mem_reg[20][27]  ( .D(n8622), .CK(CLK), .Q(net254282), .QN(
        n36777) );
  DFF_X1 \DRAM_mem_reg[20][26]  ( .D(n8621), .CK(CLK), .Q(net254281), .QN(
        n36776) );
  DFF_X1 \DRAM_mem_reg[20][25]  ( .D(n8620), .CK(CLK), .Q(net254280), .QN(
        n36775) );
  DFF_X1 \DRAM_mem_reg[20][24]  ( .D(n8619), .CK(CLK), .Q(net254279), .QN(
        n36774) );
  DFF_X1 \DRAM_mem_reg[20][23]  ( .D(n8618), .CK(CLK), .Q(net254278), .QN(
        n37069) );
  DFF_X1 \DRAM_mem_reg[20][22]  ( .D(n8617), .CK(CLK), .Q(net254277), .QN(
        n37068) );
  DFF_X1 \DRAM_mem_reg[20][21]  ( .D(n8616), .CK(CLK), .Q(net254276), .QN(
        n37067) );
  DFF_X1 \DRAM_mem_reg[20][20]  ( .D(n8615), .CK(CLK), .Q(net254275), .QN(
        n37066) );
  DFF_X1 \DRAM_mem_reg[20][19]  ( .D(n8614), .CK(CLK), .Q(net254274), .QN(
        n37065) );
  DFF_X1 \DRAM_mem_reg[20][18]  ( .D(n8613), .CK(CLK), .Q(net254273), .QN(
        n37064) );
  DFF_X1 \DRAM_mem_reg[20][17]  ( .D(n8612), .CK(CLK), .Q(net254272), .QN(
        n37063) );
  DFF_X1 \DRAM_mem_reg[20][16]  ( .D(n8611), .CK(CLK), .Q(net254271), .QN(
        n37062) );
  DFF_X1 \DRAM_mem_reg[20][15]  ( .D(n8610), .CK(CLK), .Q(net254270), .QN(
        n37061) );
  DFF_X1 \DRAM_mem_reg[20][14]  ( .D(n8609), .CK(CLK), .Q(net254269), .QN(
        n37060) );
  DFF_X1 \DRAM_mem_reg[20][13]  ( .D(n8608), .CK(CLK), .Q(net254268), .QN(
        n37059) );
  DFF_X1 \DRAM_mem_reg[20][12]  ( .D(n8607), .CK(CLK), .Q(net254267), .QN(
        n37058) );
  DFF_X1 \DRAM_mem_reg[20][11]  ( .D(n8606), .CK(CLK), .Q(net254266), .QN(
        n37057) );
  DFF_X1 \DRAM_mem_reg[20][10]  ( .D(n8605), .CK(CLK), .Q(net254265), .QN(
        n37056) );
  DFF_X1 \DRAM_mem_reg[20][9]  ( .D(n8604), .CK(CLK), .Q(net254264), .QN(
        n37055) );
  DFF_X1 \DRAM_mem_reg[20][8]  ( .D(n8603), .CK(CLK), .Q(net254263), .QN(
        n37054) );
  DFF_X1 \DRAM_mem_reg[20][7]  ( .D(n8602), .CK(CLK), .Q(net254262), .QN(
        n37053) );
  DFF_X1 \DRAM_mem_reg[20][6]  ( .D(n8601), .CK(CLK), .Q(net254261), .QN(
        n37052) );
  DFF_X1 \DRAM_mem_reg[20][5]  ( .D(n8600), .CK(CLK), .Q(net254260), .QN(
        n37051) );
  DFF_X1 \DRAM_mem_reg[20][4]  ( .D(n8599), .CK(CLK), .Q(net254259), .QN(
        n37050) );
  DFF_X1 \DRAM_mem_reg[20][3]  ( .D(n8598), .CK(CLK), .Q(net254258), .QN(
        n37049) );
  DFF_X1 \DRAM_mem_reg[20][2]  ( .D(n8597), .CK(CLK), .Q(net254257), .QN(
        n37048) );
  DFF_X1 \DRAM_mem_reg[20][1]  ( .D(n8596), .CK(CLK), .Q(net254256), .QN(
        n37047) );
  DFF_X1 \DRAM_mem_reg[20][0]  ( .D(n8595), .CK(CLK), .Q(net254255), .QN(
        n37046) );
  DFF_X1 \DRAM_mem_reg[21][31]  ( .D(n8594), .CK(CLK), .QN(n35410) );
  DFF_X1 \DRAM_mem_reg[21][30]  ( .D(n8593), .CK(CLK), .QN(n35401) );
  DFF_X1 \DRAM_mem_reg[21][29]  ( .D(n8592), .CK(CLK), .QN(n35392) );
  DFF_X1 \DRAM_mem_reg[21][28]  ( .D(n8591), .CK(CLK), .QN(n35383) );
  DFF_X1 \DRAM_mem_reg[21][27]  ( .D(n8590), .CK(CLK), .QN(n35374) );
  DFF_X1 \DRAM_mem_reg[21][26]  ( .D(n8589), .CK(CLK), .QN(n35365) );
  DFF_X1 \DRAM_mem_reg[21][25]  ( .D(n8588), .CK(CLK), .QN(n35356) );
  DFF_X1 \DRAM_mem_reg[21][24]  ( .D(n8587), .CK(CLK), .QN(n35347) );
  DFF_X1 \DRAM_mem_reg[21][23]  ( .D(n8586), .CK(CLK), .QN(n35509) );
  DFF_X1 \DRAM_mem_reg[21][22]  ( .D(n8585), .CK(CLK), .QN(n35505) );
  DFF_X1 \DRAM_mem_reg[21][21]  ( .D(n8584), .CK(CLK), .QN(n35501) );
  DFF_X1 \DRAM_mem_reg[21][20]  ( .D(n8583), .CK(CLK), .QN(n35497) );
  DFF_X1 \DRAM_mem_reg[21][19]  ( .D(n8582), .CK(CLK), .QN(n35493) );
  DFF_X1 \DRAM_mem_reg[21][18]  ( .D(n8581), .CK(CLK), .QN(n35489) );
  DFF_X1 \DRAM_mem_reg[21][17]  ( .D(n8580), .CK(CLK), .QN(n35485) );
  DFF_X1 \DRAM_mem_reg[21][16]  ( .D(n8579), .CK(CLK), .QN(n35481) );
  DFF_X1 \DRAM_mem_reg[21][15]  ( .D(n8578), .CK(CLK), .QN(n35477) );
  DFF_X1 \DRAM_mem_reg[21][14]  ( .D(n8577), .CK(CLK), .QN(n35473) );
  DFF_X1 \DRAM_mem_reg[21][13]  ( .D(n8576), .CK(CLK), .QN(n35469) );
  DFF_X1 \DRAM_mem_reg[21][12]  ( .D(n8575), .CK(CLK), .QN(n35465) );
  DFF_X1 \DRAM_mem_reg[21][11]  ( .D(n8574), .CK(CLK), .QN(n35461) );
  DFF_X1 \DRAM_mem_reg[21][10]  ( .D(n8573), .CK(CLK), .QN(n35457) );
  DFF_X1 \DRAM_mem_reg[21][9]  ( .D(n8572), .CK(CLK), .QN(n35453) );
  DFF_X1 \DRAM_mem_reg[21][8]  ( .D(n8571), .CK(CLK), .QN(n35449) );
  DFF_X1 \DRAM_mem_reg[21][7]  ( .D(n8570), .CK(CLK), .QN(n35445) );
  DFF_X1 \DRAM_mem_reg[21][6]  ( .D(n8569), .CK(CLK), .QN(n35441) );
  DFF_X1 \DRAM_mem_reg[21][5]  ( .D(n8568), .CK(CLK), .QN(n35437) );
  DFF_X1 \DRAM_mem_reg[21][4]  ( .D(n8567), .CK(CLK), .QN(n35433) );
  DFF_X1 \DRAM_mem_reg[21][3]  ( .D(n8566), .CK(CLK), .QN(n35429) );
  DFF_X1 \DRAM_mem_reg[21][2]  ( .D(n8565), .CK(CLK), .QN(n35425) );
  DFF_X1 \DRAM_mem_reg[21][1]  ( .D(n8564), .CK(CLK), .QN(n35421) );
  DFF_X1 \DRAM_mem_reg[21][0]  ( .D(n8563), .CK(CLK), .QN(n35417) );
  DFF_X1 \DRAM_mem_reg[22][31]  ( .D(n8562), .CK(CLK), .QN(n35925) );
  DFF_X1 \DRAM_mem_reg[22][30]  ( .D(n8561), .CK(CLK), .QN(n35916) );
  DFF_X1 \DRAM_mem_reg[22][29]  ( .D(n8560), .CK(CLK), .QN(n35907) );
  DFF_X1 \DRAM_mem_reg[22][28]  ( .D(n8559), .CK(CLK), .QN(n35898) );
  DFF_X1 \DRAM_mem_reg[22][27]  ( .D(n8558), .CK(CLK), .QN(n35889) );
  DFF_X1 \DRAM_mem_reg[22][26]  ( .D(n8557), .CK(CLK), .QN(n35880) );
  DFF_X1 \DRAM_mem_reg[22][25]  ( .D(n8556), .CK(CLK), .QN(n35871) );
  DFF_X1 \DRAM_mem_reg[22][24]  ( .D(n8555), .CK(CLK), .QN(n35862) );
  DFF_X1 \DRAM_mem_reg[22][23]  ( .D(n8554), .CK(CLK), .QN(n36173) );
  DFF_X1 \DRAM_mem_reg[22][22]  ( .D(n8553), .CK(CLK), .QN(n36171) );
  DFF_X1 \DRAM_mem_reg[22][21]  ( .D(n8552), .CK(CLK), .QN(n36169) );
  DFF_X1 \DRAM_mem_reg[22][20]  ( .D(n8551), .CK(CLK), .QN(n36167) );
  DFF_X1 \DRAM_mem_reg[22][19]  ( .D(n8550), .CK(CLK), .QN(n36165) );
  DFF_X1 \DRAM_mem_reg[22][18]  ( .D(n8549), .CK(CLK), .QN(n36163) );
  DFF_X1 \DRAM_mem_reg[22][17]  ( .D(n8548), .CK(CLK), .QN(n36161) );
  DFF_X1 \DRAM_mem_reg[22][16]  ( .D(n8547), .CK(CLK), .QN(n36159) );
  DFF_X1 \DRAM_mem_reg[22][15]  ( .D(n8546), .CK(CLK), .QN(n36157) );
  DFF_X1 \DRAM_mem_reg[22][14]  ( .D(n8545), .CK(CLK), .QN(n36155) );
  DFF_X1 \DRAM_mem_reg[22][13]  ( .D(n8544), .CK(CLK), .QN(n36153) );
  DFF_X1 \DRAM_mem_reg[22][12]  ( .D(n8543), .CK(CLK), .QN(n36151) );
  DFF_X1 \DRAM_mem_reg[22][11]  ( .D(n8542), .CK(CLK), .QN(n36149) );
  DFF_X1 \DRAM_mem_reg[22][10]  ( .D(n8541), .CK(CLK), .QN(n36147) );
  DFF_X1 \DRAM_mem_reg[22][9]  ( .D(n8540), .CK(CLK), .QN(n36145) );
  DFF_X1 \DRAM_mem_reg[22][8]  ( .D(n8539), .CK(CLK), .QN(n36143) );
  DFF_X1 \DRAM_mem_reg[22][7]  ( .D(n8538), .CK(CLK), .QN(n36141) );
  DFF_X1 \DRAM_mem_reg[22][6]  ( .D(n8537), .CK(CLK), .QN(n36139) );
  DFF_X1 \DRAM_mem_reg[22][5]  ( .D(n8536), .CK(CLK), .QN(n36137) );
  DFF_X1 \DRAM_mem_reg[22][4]  ( .D(n8535), .CK(CLK), .QN(n36135) );
  DFF_X1 \DRAM_mem_reg[22][3]  ( .D(n8534), .CK(CLK), .QN(n36133) );
  DFF_X1 \DRAM_mem_reg[22][2]  ( .D(n8533), .CK(CLK), .QN(n36131) );
  DFF_X1 \DRAM_mem_reg[22][1]  ( .D(n8532), .CK(CLK), .QN(n36129) );
  DFF_X1 \DRAM_mem_reg[22][0]  ( .D(n8531), .CK(CLK), .QN(n36127) );
  DFF_X1 \DRAM_mem_reg[23][31]  ( .D(n8530), .CK(CLK), .Q(net254254), .QN(
        n37157) );
  DFF_X1 \DRAM_mem_reg[23][30]  ( .D(n8529), .CK(CLK), .Q(net254253), .QN(
        n37156) );
  DFF_X1 \DRAM_mem_reg[23][29]  ( .D(n8528), .CK(CLK), .Q(net254252), .QN(
        n37155) );
  DFF_X1 \DRAM_mem_reg[23][28]  ( .D(n8527), .CK(CLK), .Q(net254251), .QN(
        n37154) );
  DFF_X1 \DRAM_mem_reg[23][27]  ( .D(n8526), .CK(CLK), .Q(net254250), .QN(
        n37153) );
  DFF_X1 \DRAM_mem_reg[23][26]  ( .D(n8525), .CK(CLK), .Q(net254249), .QN(
        n37152) );
  DFF_X1 \DRAM_mem_reg[23][25]  ( .D(n8524), .CK(CLK), .Q(net254248), .QN(
        n37151) );
  DFF_X1 \DRAM_mem_reg[23][24]  ( .D(n8523), .CK(CLK), .Q(net254247), .QN(
        n37150) );
  DFF_X1 \DRAM_mem_reg[23][23]  ( .D(n8522), .CK(CLK), .Q(net254246), .QN(
        n37429) );
  DFF_X1 \DRAM_mem_reg[23][22]  ( .D(n8521), .CK(CLK), .Q(net254245), .QN(
        n37428) );
  DFF_X1 \DRAM_mem_reg[23][21]  ( .D(n8520), .CK(CLK), .Q(net254244), .QN(
        n37427) );
  DFF_X1 \DRAM_mem_reg[23][20]  ( .D(n8519), .CK(CLK), .Q(net254243), .QN(
        n37426) );
  DFF_X1 \DRAM_mem_reg[23][19]  ( .D(n8518), .CK(CLK), .Q(net254242), .QN(
        n37425) );
  DFF_X1 \DRAM_mem_reg[23][18]  ( .D(n8517), .CK(CLK), .Q(net254241), .QN(
        n37424) );
  DFF_X1 \DRAM_mem_reg[23][17]  ( .D(n8516), .CK(CLK), .Q(net254240), .QN(
        n37423) );
  DFF_X1 \DRAM_mem_reg[23][16]  ( .D(n8515), .CK(CLK), .Q(net254239), .QN(
        n37422) );
  DFF_X1 \DRAM_mem_reg[23][15]  ( .D(n8514), .CK(CLK), .Q(net254238), .QN(
        n37421) );
  DFF_X1 \DRAM_mem_reg[23][14]  ( .D(n8513), .CK(CLK), .Q(net254237), .QN(
        n37420) );
  DFF_X1 \DRAM_mem_reg[23][13]  ( .D(n8512), .CK(CLK), .Q(net254236), .QN(
        n37419) );
  DFF_X1 \DRAM_mem_reg[23][12]  ( .D(n8511), .CK(CLK), .Q(net254235), .QN(
        n37418) );
  DFF_X1 \DRAM_mem_reg[23][11]  ( .D(n8510), .CK(CLK), .Q(net254234), .QN(
        n37417) );
  DFF_X1 \DRAM_mem_reg[23][10]  ( .D(n8509), .CK(CLK), .Q(net254233), .QN(
        n37416) );
  DFF_X1 \DRAM_mem_reg[23][9]  ( .D(n8508), .CK(CLK), .Q(net254232), .QN(
        n37415) );
  DFF_X1 \DRAM_mem_reg[23][8]  ( .D(n8507), .CK(CLK), .Q(net254231), .QN(
        n37414) );
  DFF_X1 \DRAM_mem_reg[23][7]  ( .D(n8506), .CK(CLK), .Q(net254230), .QN(
        n37413) );
  DFF_X1 \DRAM_mem_reg[23][6]  ( .D(n8505), .CK(CLK), .Q(net254229), .QN(
        n37412) );
  DFF_X1 \DRAM_mem_reg[23][5]  ( .D(n8504), .CK(CLK), .Q(net254228), .QN(
        n37411) );
  DFF_X1 \DRAM_mem_reg[23][4]  ( .D(n8503), .CK(CLK), .Q(net254227), .QN(
        n37410) );
  DFF_X1 \DRAM_mem_reg[23][3]  ( .D(n8502), .CK(CLK), .Q(net254226), .QN(
        n37409) );
  DFF_X1 \DRAM_mem_reg[23][2]  ( .D(n8501), .CK(CLK), .Q(net254225), .QN(
        n37408) );
  DFF_X1 \DRAM_mem_reg[23][1]  ( .D(n8500), .CK(CLK), .Q(net254224), .QN(
        n37407) );
  DFF_X1 \DRAM_mem_reg[23][0]  ( .D(n8499), .CK(CLK), .Q(net254223), .QN(
        n37406) );
  DFF_X1 \DRAM_mem_reg[24][31]  ( .D(n8498), .CK(CLK), .QN(n36436) );
  DFF_X1 \DRAM_mem_reg[24][30]  ( .D(n8497), .CK(CLK), .QN(n36427) );
  DFF_X1 \DRAM_mem_reg[24][29]  ( .D(n8496), .CK(CLK), .QN(n36418) );
  DFF_X1 \DRAM_mem_reg[24][28]  ( .D(n8495), .CK(CLK), .QN(n36409) );
  DFF_X1 \DRAM_mem_reg[24][27]  ( .D(n8494), .CK(CLK), .QN(n36400) );
  DFF_X1 \DRAM_mem_reg[24][26]  ( .D(n8493), .CK(CLK), .QN(n36391) );
  DFF_X1 \DRAM_mem_reg[24][25]  ( .D(n8492), .CK(CLK), .QN(n36382) );
  DFF_X1 \DRAM_mem_reg[24][24]  ( .D(n8491), .CK(CLK), .QN(n36373) );
  DFF_X1 \DRAM_mem_reg[24][23]  ( .D(n8490), .CK(CLK), .QN(n36637) );
  DFF_X1 \DRAM_mem_reg[24][22]  ( .D(n8489), .CK(CLK), .QN(n36635) );
  DFF_X1 \DRAM_mem_reg[24][21]  ( .D(n8488), .CK(CLK), .QN(n36633) );
  DFF_X1 \DRAM_mem_reg[24][20]  ( .D(n8487), .CK(CLK), .QN(n36631) );
  DFF_X1 \DRAM_mem_reg[24][19]  ( .D(n8486), .CK(CLK), .QN(n36629) );
  DFF_X1 \DRAM_mem_reg[24][18]  ( .D(n8485), .CK(CLK), .QN(n36627) );
  DFF_X1 \DRAM_mem_reg[24][17]  ( .D(n8484), .CK(CLK), .QN(n36625) );
  DFF_X1 \DRAM_mem_reg[24][16]  ( .D(n8483), .CK(CLK), .QN(n36623) );
  DFF_X1 \DRAM_mem_reg[24][15]  ( .D(n8482), .CK(CLK), .QN(n36621) );
  DFF_X1 \DRAM_mem_reg[24][14]  ( .D(n8481), .CK(CLK), .QN(n36619) );
  DFF_X1 \DRAM_mem_reg[24][13]  ( .D(n8480), .CK(CLK), .QN(n36617) );
  DFF_X1 \DRAM_mem_reg[24][12]  ( .D(n8479), .CK(CLK), .QN(n36615) );
  DFF_X1 \DRAM_mem_reg[24][11]  ( .D(n8478), .CK(CLK), .QN(n36613) );
  DFF_X1 \DRAM_mem_reg[24][10]  ( .D(n8477), .CK(CLK), .QN(n36611) );
  DFF_X1 \DRAM_mem_reg[24][9]  ( .D(n8476), .CK(CLK), .QN(n36609) );
  DFF_X1 \DRAM_mem_reg[24][8]  ( .D(n8475), .CK(CLK), .QN(n36607) );
  DFF_X1 \DRAM_mem_reg[24][7]  ( .D(n8474), .CK(CLK), .QN(n36605) );
  DFF_X1 \DRAM_mem_reg[24][6]  ( .D(n8473), .CK(CLK), .QN(n36603) );
  DFF_X1 \DRAM_mem_reg[24][5]  ( .D(n8472), .CK(CLK), .QN(n36601) );
  DFF_X1 \DRAM_mem_reg[24][4]  ( .D(n8471), .CK(CLK), .QN(n36599) );
  DFF_X1 \DRAM_mem_reg[24][3]  ( .D(n8470), .CK(CLK), .QN(n36597) );
  DFF_X1 \DRAM_mem_reg[24][2]  ( .D(n8469), .CK(CLK), .QN(n36595) );
  DFF_X1 \DRAM_mem_reg[24][1]  ( .D(n8468), .CK(CLK), .QN(n36593) );
  DFF_X1 \DRAM_mem_reg[24][0]  ( .D(n8467), .CK(CLK), .QN(n36591) );
  DFF_X1 \DRAM_mem_reg[25][31]  ( .D(n8466), .CK(CLK), .Q(net254222), .QN(
        n36773) );
  DFF_X1 \DRAM_mem_reg[25][30]  ( .D(n8465), .CK(CLK), .Q(net254221), .QN(
        n36772) );
  DFF_X1 \DRAM_mem_reg[25][29]  ( .D(n8464), .CK(CLK), .Q(net254220), .QN(
        n36771) );
  DFF_X1 \DRAM_mem_reg[25][28]  ( .D(n8463), .CK(CLK), .Q(net254219), .QN(
        n36770) );
  DFF_X1 \DRAM_mem_reg[25][27]  ( .D(n8462), .CK(CLK), .Q(net254218), .QN(
        n36769) );
  DFF_X1 \DRAM_mem_reg[25][26]  ( .D(n8461), .CK(CLK), .Q(net254217), .QN(
        n36768) );
  DFF_X1 \DRAM_mem_reg[25][25]  ( .D(n8460), .CK(CLK), .Q(net254216), .QN(
        n36767) );
  DFF_X1 \DRAM_mem_reg[25][24]  ( .D(n8459), .CK(CLK), .Q(net254215), .QN(
        n36766) );
  DFF_X1 \DRAM_mem_reg[25][23]  ( .D(n8458), .CK(CLK), .Q(net254214), .QN(
        n37045) );
  DFF_X1 \DRAM_mem_reg[25][22]  ( .D(n8457), .CK(CLK), .Q(net254213), .QN(
        n37044) );
  DFF_X1 \DRAM_mem_reg[25][21]  ( .D(n8456), .CK(CLK), .Q(net254212), .QN(
        n37043) );
  DFF_X1 \DRAM_mem_reg[25][20]  ( .D(n8455), .CK(CLK), .Q(net254211), .QN(
        n37042) );
  DFF_X1 \DRAM_mem_reg[25][19]  ( .D(n8454), .CK(CLK), .Q(net254210), .QN(
        n37041) );
  DFF_X1 \DRAM_mem_reg[25][18]  ( .D(n8453), .CK(CLK), .Q(net254209), .QN(
        n37040) );
  DFF_X1 \DRAM_mem_reg[25][17]  ( .D(n8452), .CK(CLK), .Q(net254208), .QN(
        n37039) );
  DFF_X1 \DRAM_mem_reg[25][16]  ( .D(n8451), .CK(CLK), .Q(net254207), .QN(
        n37038) );
  DFF_X1 \DRAM_mem_reg[25][15]  ( .D(n8450), .CK(CLK), .Q(net254206), .QN(
        n37037) );
  DFF_X1 \DRAM_mem_reg[25][14]  ( .D(n8449), .CK(CLK), .Q(net254205), .QN(
        n37036) );
  DFF_X1 \DRAM_mem_reg[25][13]  ( .D(n8448), .CK(CLK), .Q(net254204), .QN(
        n37035) );
  DFF_X1 \DRAM_mem_reg[25][12]  ( .D(n8447), .CK(CLK), .Q(net254203), .QN(
        n37034) );
  DFF_X1 \DRAM_mem_reg[25][11]  ( .D(n8446), .CK(CLK), .Q(net254202), .QN(
        n37033) );
  DFF_X1 \DRAM_mem_reg[25][10]  ( .D(n8445), .CK(CLK), .Q(net254201), .QN(
        n37032) );
  DFF_X1 \DRAM_mem_reg[25][9]  ( .D(n8444), .CK(CLK), .Q(net254200), .QN(
        n37031) );
  DFF_X1 \DRAM_mem_reg[25][8]  ( .D(n8443), .CK(CLK), .Q(net254199), .QN(
        n37030) );
  DFF_X1 \DRAM_mem_reg[25][7]  ( .D(n8442), .CK(CLK), .Q(net254198), .QN(
        n37029) );
  DFF_X1 \DRAM_mem_reg[25][6]  ( .D(n8441), .CK(CLK), .Q(net254197), .QN(
        n37028) );
  DFF_X1 \DRAM_mem_reg[25][5]  ( .D(n8440), .CK(CLK), .Q(net254196), .QN(
        n37027) );
  DFF_X1 \DRAM_mem_reg[25][4]  ( .D(n8439), .CK(CLK), .Q(net254195), .QN(
        n37026) );
  DFF_X1 \DRAM_mem_reg[25][3]  ( .D(n8438), .CK(CLK), .Q(net254194), .QN(
        n37025) );
  DFF_X1 \DRAM_mem_reg[25][2]  ( .D(n8437), .CK(CLK), .Q(net254193), .QN(
        n37024) );
  DFF_X1 \DRAM_mem_reg[25][1]  ( .D(n8436), .CK(CLK), .Q(net254192), .QN(
        n37023) );
  DFF_X1 \DRAM_mem_reg[25][0]  ( .D(n8435), .CK(CLK), .Q(net254191), .QN(
        n37022) );
  DFF_X1 \DRAM_mem_reg[26][31]  ( .D(n8434), .CK(CLK), .QN(n35407) );
  DFF_X1 \DRAM_mem_reg[26][30]  ( .D(n8433), .CK(CLK), .QN(n35398) );
  DFF_X1 \DRAM_mem_reg[26][29]  ( .D(n8432), .CK(CLK), .QN(n35389) );
  DFF_X1 \DRAM_mem_reg[26][28]  ( .D(n8431), .CK(CLK), .QN(n35380) );
  DFF_X1 \DRAM_mem_reg[26][27]  ( .D(n8430), .CK(CLK), .QN(n35371) );
  DFF_X1 \DRAM_mem_reg[26][26]  ( .D(n8429), .CK(CLK), .QN(n35362) );
  DFF_X1 \DRAM_mem_reg[26][25]  ( .D(n8428), .CK(CLK), .QN(n35353) );
  DFF_X1 \DRAM_mem_reg[26][24]  ( .D(n8427), .CK(CLK), .QN(n35344) );
  DFF_X1 \DRAM_mem_reg[26][23]  ( .D(n8426), .CK(CLK), .QN(n35564) );
  DFF_X1 \DRAM_mem_reg[26][22]  ( .D(n8425), .CK(CLK), .QN(n35562) );
  DFF_X1 \DRAM_mem_reg[26][21]  ( .D(n8424), .CK(CLK), .QN(n35560) );
  DFF_X1 \DRAM_mem_reg[26][20]  ( .D(n8423), .CK(CLK), .QN(n35558) );
  DFF_X1 \DRAM_mem_reg[26][19]  ( .D(n8422), .CK(CLK), .QN(n35556) );
  DFF_X1 \DRAM_mem_reg[26][18]  ( .D(n8421), .CK(CLK), .QN(n35554) );
  DFF_X1 \DRAM_mem_reg[26][17]  ( .D(n8420), .CK(CLK), .QN(n35552) );
  DFF_X1 \DRAM_mem_reg[26][16]  ( .D(n8419), .CK(CLK), .QN(n35550) );
  DFF_X1 \DRAM_mem_reg[26][15]  ( .D(n8418), .CK(CLK), .QN(n35548) );
  DFF_X1 \DRAM_mem_reg[26][14]  ( .D(n8417), .CK(CLK), .QN(n35546) );
  DFF_X1 \DRAM_mem_reg[26][13]  ( .D(n8416), .CK(CLK), .QN(n35544) );
  DFF_X1 \DRAM_mem_reg[26][12]  ( .D(n8415), .CK(CLK), .QN(n35542) );
  DFF_X1 \DRAM_mem_reg[26][11]  ( .D(n8414), .CK(CLK), .QN(n35540) );
  DFF_X1 \DRAM_mem_reg[26][10]  ( .D(n8413), .CK(CLK), .QN(n35538) );
  DFF_X1 \DRAM_mem_reg[26][9]  ( .D(n8412), .CK(CLK), .QN(n35536) );
  DFF_X1 \DRAM_mem_reg[26][8]  ( .D(n8411), .CK(CLK), .QN(n35534) );
  DFF_X1 \DRAM_mem_reg[26][7]  ( .D(n8410), .CK(CLK), .QN(n35532) );
  DFF_X1 \DRAM_mem_reg[26][6]  ( .D(n8409), .CK(CLK), .QN(n35530) );
  DFF_X1 \DRAM_mem_reg[26][5]  ( .D(n8408), .CK(CLK), .QN(n35528) );
  DFF_X1 \DRAM_mem_reg[26][4]  ( .D(n8407), .CK(CLK), .QN(n35526) );
  DFF_X1 \DRAM_mem_reg[26][3]  ( .D(n8406), .CK(CLK), .QN(n35524) );
  DFF_X1 \DRAM_mem_reg[26][2]  ( .D(n8405), .CK(CLK), .QN(n35522) );
  DFF_X1 \DRAM_mem_reg[26][1]  ( .D(n8404), .CK(CLK), .QN(n35520) );
  DFF_X1 \DRAM_mem_reg[26][0]  ( .D(n8403), .CK(CLK), .QN(n35518) );
  DFF_X1 \DRAM_mem_reg[27][31]  ( .D(n8402), .CK(CLK), .QN(n35918) );
  DFF_X1 \DRAM_mem_reg[27][30]  ( .D(n8401), .CK(CLK), .QN(n35909) );
  DFF_X1 \DRAM_mem_reg[27][29]  ( .D(n8400), .CK(CLK), .QN(n35900) );
  DFF_X1 \DRAM_mem_reg[27][28]  ( .D(n8399), .CK(CLK), .QN(n35891) );
  DFF_X1 \DRAM_mem_reg[27][27]  ( .D(n8398), .CK(CLK), .QN(n35882) );
  DFF_X1 \DRAM_mem_reg[27][26]  ( .D(n8397), .CK(CLK), .QN(n35873) );
  DFF_X1 \DRAM_mem_reg[27][25]  ( .D(n8396), .CK(CLK), .QN(n35864) );
  DFF_X1 \DRAM_mem_reg[27][24]  ( .D(n8395), .CK(CLK), .QN(n35855) );
  DFF_X1 \DRAM_mem_reg[27][23]  ( .D(n8394), .CK(CLK), .QN(n36020) );
  DFF_X1 \DRAM_mem_reg[27][22]  ( .D(n8393), .CK(CLK), .QN(n36016) );
  DFF_X1 \DRAM_mem_reg[27][21]  ( .D(n8392), .CK(CLK), .QN(n36012) );
  DFF_X1 \DRAM_mem_reg[27][20]  ( .D(n8391), .CK(CLK), .QN(n36008) );
  DFF_X1 \DRAM_mem_reg[27][19]  ( .D(n8390), .CK(CLK), .QN(n36004) );
  DFF_X1 \DRAM_mem_reg[27][18]  ( .D(n8389), .CK(CLK), .QN(n36000) );
  DFF_X1 \DRAM_mem_reg[27][17]  ( .D(n8388), .CK(CLK), .QN(n35996) );
  DFF_X1 \DRAM_mem_reg[27][16]  ( .D(n8387), .CK(CLK), .QN(n35992) );
  DFF_X1 \DRAM_mem_reg[27][15]  ( .D(n8386), .CK(CLK), .QN(n35988) );
  DFF_X1 \DRAM_mem_reg[27][14]  ( .D(n8385), .CK(CLK), .QN(n35984) );
  DFF_X1 \DRAM_mem_reg[27][13]  ( .D(n8384), .CK(CLK), .QN(n35980) );
  DFF_X1 \DRAM_mem_reg[27][12]  ( .D(n8383), .CK(CLK), .QN(n35976) );
  DFF_X1 \DRAM_mem_reg[27][11]  ( .D(n8382), .CK(CLK), .QN(n35972) );
  DFF_X1 \DRAM_mem_reg[27][10]  ( .D(n8381), .CK(CLK), .QN(n35968) );
  DFF_X1 \DRAM_mem_reg[27][9]  ( .D(n8380), .CK(CLK), .QN(n35964) );
  DFF_X1 \DRAM_mem_reg[27][8]  ( .D(n8379), .CK(CLK), .QN(n35960) );
  DFF_X1 \DRAM_mem_reg[27][7]  ( .D(n8378), .CK(CLK), .QN(n35956) );
  DFF_X1 \DRAM_mem_reg[27][6]  ( .D(n8377), .CK(CLK), .QN(n35952) );
  DFF_X1 \DRAM_mem_reg[27][5]  ( .D(n8376), .CK(CLK), .QN(n35948) );
  DFF_X1 \DRAM_mem_reg[27][4]  ( .D(n8375), .CK(CLK), .QN(n35944) );
  DFF_X1 \DRAM_mem_reg[27][3]  ( .D(n8374), .CK(CLK), .QN(n35940) );
  DFF_X1 \DRAM_mem_reg[27][2]  ( .D(n8373), .CK(CLK), .QN(n35936) );
  DFF_X1 \DRAM_mem_reg[27][1]  ( .D(n8372), .CK(CLK), .QN(n35932) );
  DFF_X1 \DRAM_mem_reg[27][0]  ( .D(n8371), .CK(CLK), .QN(n35928) );
  DFF_X1 \DRAM_mem_reg[28][31]  ( .D(n8370), .CK(CLK), .Q(net254190), .QN(
        n37149) );
  DFF_X1 \DRAM_mem_reg[28][30]  ( .D(n8369), .CK(CLK), .Q(net254189), .QN(
        n37148) );
  DFF_X1 \DRAM_mem_reg[28][29]  ( .D(n8368), .CK(CLK), .Q(net254188), .QN(
        n37147) );
  DFF_X1 \DRAM_mem_reg[28][28]  ( .D(n8367), .CK(CLK), .Q(net254187), .QN(
        n37146) );
  DFF_X1 \DRAM_mem_reg[28][27]  ( .D(n8366), .CK(CLK), .Q(net254186), .QN(
        n37145) );
  DFF_X1 \DRAM_mem_reg[28][26]  ( .D(n8365), .CK(CLK), .Q(net254185), .QN(
        n37144) );
  DFF_X1 \DRAM_mem_reg[28][25]  ( .D(n8364), .CK(CLK), .Q(net254184), .QN(
        n37143) );
  DFF_X1 \DRAM_mem_reg[28][24]  ( .D(n8363), .CK(CLK), .Q(net254183), .QN(
        n37142) );
  DFF_X1 \DRAM_mem_reg[28][23]  ( .D(n8362), .CK(CLK), .Q(net254182), .QN(
        n37405) );
  DFF_X1 \DRAM_mem_reg[28][22]  ( .D(n8361), .CK(CLK), .Q(net254181), .QN(
        n37404) );
  DFF_X1 \DRAM_mem_reg[28][21]  ( .D(n8360), .CK(CLK), .Q(net254180), .QN(
        n37403) );
  DFF_X1 \DRAM_mem_reg[28][20]  ( .D(n8359), .CK(CLK), .Q(net254179), .QN(
        n37402) );
  DFF_X1 \DRAM_mem_reg[28][19]  ( .D(n8358), .CK(CLK), .Q(net254178), .QN(
        n37401) );
  DFF_X1 \DRAM_mem_reg[28][18]  ( .D(n8357), .CK(CLK), .Q(net254177), .QN(
        n37400) );
  DFF_X1 \DRAM_mem_reg[28][17]  ( .D(n8356), .CK(CLK), .Q(net254176), .QN(
        n37399) );
  DFF_X1 \DRAM_mem_reg[28][16]  ( .D(n8355), .CK(CLK), .Q(net254175), .QN(
        n37398) );
  DFF_X1 \DRAM_mem_reg[28][15]  ( .D(n8354), .CK(CLK), .Q(net254174), .QN(
        n37397) );
  DFF_X1 \DRAM_mem_reg[28][14]  ( .D(n8353), .CK(CLK), .Q(net254173), .QN(
        n37396) );
  DFF_X1 \DRAM_mem_reg[28][13]  ( .D(n8352), .CK(CLK), .Q(net254172), .QN(
        n37395) );
  DFF_X1 \DRAM_mem_reg[28][12]  ( .D(n8351), .CK(CLK), .Q(net254171), .QN(
        n37394) );
  DFF_X1 \DRAM_mem_reg[28][11]  ( .D(n8350), .CK(CLK), .Q(net254170), .QN(
        n37393) );
  DFF_X1 \DRAM_mem_reg[28][10]  ( .D(n8349), .CK(CLK), .Q(net254169), .QN(
        n37392) );
  DFF_X1 \DRAM_mem_reg[28][9]  ( .D(n8348), .CK(CLK), .Q(net254168), .QN(
        n37391) );
  DFF_X1 \DRAM_mem_reg[28][8]  ( .D(n8347), .CK(CLK), .Q(net254167), .QN(
        n37390) );
  DFF_X1 \DRAM_mem_reg[28][7]  ( .D(n8346), .CK(CLK), .Q(net254166), .QN(
        n37389) );
  DFF_X1 \DRAM_mem_reg[28][6]  ( .D(n8345), .CK(CLK), .Q(net254165), .QN(
        n37388) );
  DFF_X1 \DRAM_mem_reg[28][5]  ( .D(n8344), .CK(CLK), .Q(net254164), .QN(
        n37387) );
  DFF_X1 \DRAM_mem_reg[28][4]  ( .D(n8343), .CK(CLK), .Q(net254163), .QN(
        n37386) );
  DFF_X1 \DRAM_mem_reg[28][3]  ( .D(n8342), .CK(CLK), .Q(net254162), .QN(
        n37385) );
  DFF_X1 \DRAM_mem_reg[28][2]  ( .D(n8341), .CK(CLK), .Q(net254161), .QN(
        n37384) );
  DFF_X1 \DRAM_mem_reg[28][1]  ( .D(n8340), .CK(CLK), .Q(net254160), .QN(
        n37383) );
  DFF_X1 \DRAM_mem_reg[28][0]  ( .D(n8339), .CK(CLK), .Q(net254159), .QN(
        n37382) );
  DFF_X1 \DRAM_mem_reg[29][31]  ( .D(n8338), .CK(CLK), .QN(n36433) );
  DFF_X1 \DRAM_mem_reg[29][30]  ( .D(n8337), .CK(CLK), .QN(n36424) );
  DFF_X1 \DRAM_mem_reg[29][29]  ( .D(n8336), .CK(CLK), .QN(n36415) );
  DFF_X1 \DRAM_mem_reg[29][28]  ( .D(n8335), .CK(CLK), .QN(n36406) );
  DFF_X1 \DRAM_mem_reg[29][27]  ( .D(n8334), .CK(CLK), .QN(n36397) );
  DFF_X1 \DRAM_mem_reg[29][26]  ( .D(n8333), .CK(CLK), .QN(n36388) );
  DFF_X1 \DRAM_mem_reg[29][25]  ( .D(n8332), .CK(CLK), .QN(n36379) );
  DFF_X1 \DRAM_mem_reg[29][24]  ( .D(n8331), .CK(CLK), .QN(n36370) );
  DFF_X1 \DRAM_mem_reg[29][23]  ( .D(n8330), .CK(CLK), .QN(n36684) );
  DFF_X1 \DRAM_mem_reg[29][22]  ( .D(n8329), .CK(CLK), .QN(n36682) );
  DFF_X1 \DRAM_mem_reg[29][21]  ( .D(n8328), .CK(CLK), .QN(n36680) );
  DFF_X1 \DRAM_mem_reg[29][20]  ( .D(n8327), .CK(CLK), .QN(n36678) );
  DFF_X1 \DRAM_mem_reg[29][19]  ( .D(n8326), .CK(CLK), .QN(n36676) );
  DFF_X1 \DRAM_mem_reg[29][18]  ( .D(n8325), .CK(CLK), .QN(n36674) );
  DFF_X1 \DRAM_mem_reg[29][17]  ( .D(n8324), .CK(CLK), .QN(n36672) );
  DFF_X1 \DRAM_mem_reg[29][16]  ( .D(n8323), .CK(CLK), .QN(n36670) );
  DFF_X1 \DRAM_mem_reg[29][15]  ( .D(n8322), .CK(CLK), .QN(n36668) );
  DFF_X1 \DRAM_mem_reg[29][14]  ( .D(n8321), .CK(CLK), .QN(n36666) );
  DFF_X1 \DRAM_mem_reg[29][13]  ( .D(n8320), .CK(CLK), .QN(n36664) );
  DFF_X1 \DRAM_mem_reg[29][12]  ( .D(n8319), .CK(CLK), .QN(n36662) );
  DFF_X1 \DRAM_mem_reg[29][11]  ( .D(n8318), .CK(CLK), .QN(n36660) );
  DFF_X1 \DRAM_mem_reg[29][10]  ( .D(n8317), .CK(CLK), .QN(n36658) );
  DFF_X1 \DRAM_mem_reg[29][9]  ( .D(n8316), .CK(CLK), .QN(n36656) );
  DFF_X1 \DRAM_mem_reg[29][8]  ( .D(n8315), .CK(CLK), .QN(n36654) );
  DFF_X1 \DRAM_mem_reg[29][7]  ( .D(n8314), .CK(CLK), .QN(n36652) );
  DFF_X1 \DRAM_mem_reg[29][6]  ( .D(n8313), .CK(CLK), .QN(n36650) );
  DFF_X1 \DRAM_mem_reg[29][5]  ( .D(n8312), .CK(CLK), .QN(n36648) );
  DFF_X1 \DRAM_mem_reg[29][4]  ( .D(n8311), .CK(CLK), .QN(n36646) );
  DFF_X1 \DRAM_mem_reg[29][3]  ( .D(n8310), .CK(CLK), .QN(n36644) );
  DFF_X1 \DRAM_mem_reg[29][2]  ( .D(n8309), .CK(CLK), .QN(n36642) );
  DFF_X1 \DRAM_mem_reg[29][1]  ( .D(n8308), .CK(CLK), .QN(n36640) );
  DFF_X1 \DRAM_mem_reg[29][0]  ( .D(n8307), .CK(CLK), .QN(n36638) );
  DFF_X1 \DRAM_mem_reg[30][31]  ( .D(n8306), .CK(CLK), .Q(net254158), .QN(
        n36765) );
  DFF_X1 \DRAM_mem_reg[30][30]  ( .D(n8305), .CK(CLK), .Q(net254157), .QN(
        n36764) );
  DFF_X1 \DRAM_mem_reg[30][29]  ( .D(n8304), .CK(CLK), .Q(net254156), .QN(
        n36763) );
  DFF_X1 \DRAM_mem_reg[30][28]  ( .D(n8303), .CK(CLK), .Q(net254155), .QN(
        n36762) );
  DFF_X1 \DRAM_mem_reg[30][27]  ( .D(n8302), .CK(CLK), .Q(net254154), .QN(
        n36761) );
  DFF_X1 \DRAM_mem_reg[30][26]  ( .D(n8301), .CK(CLK), .Q(net254153), .QN(
        n36760) );
  DFF_X1 \DRAM_mem_reg[30][25]  ( .D(n8300), .CK(CLK), .Q(net254152), .QN(
        n36759) );
  DFF_X1 \DRAM_mem_reg[30][24]  ( .D(n8299), .CK(CLK), .Q(net254151), .QN(
        n36758) );
  DFF_X1 \DRAM_mem_reg[30][23]  ( .D(n8298), .CK(CLK), .Q(net254150), .QN(
        n37021) );
  DFF_X1 \DRAM_mem_reg[30][22]  ( .D(n8297), .CK(CLK), .Q(net254149), .QN(
        n37020) );
  DFF_X1 \DRAM_mem_reg[30][21]  ( .D(n8296), .CK(CLK), .Q(net254148), .QN(
        n37019) );
  DFF_X1 \DRAM_mem_reg[30][20]  ( .D(n8295), .CK(CLK), .Q(net254147), .QN(
        n37018) );
  DFF_X1 \DRAM_mem_reg[30][19]  ( .D(n8294), .CK(CLK), .Q(net254146), .QN(
        n37017) );
  DFF_X1 \DRAM_mem_reg[30][18]  ( .D(n8293), .CK(CLK), .Q(net254145), .QN(
        n37016) );
  DFF_X1 \DRAM_mem_reg[30][17]  ( .D(n8292), .CK(CLK), .Q(net254144), .QN(
        n37015) );
  DFF_X1 \DRAM_mem_reg[30][16]  ( .D(n8291), .CK(CLK), .Q(net254143), .QN(
        n37014) );
  DFF_X1 \DRAM_mem_reg[30][15]  ( .D(n8290), .CK(CLK), .Q(net254142), .QN(
        n37013) );
  DFF_X1 \DRAM_mem_reg[30][14]  ( .D(n8289), .CK(CLK), .Q(net254141), .QN(
        n37012) );
  DFF_X1 \DRAM_mem_reg[30][13]  ( .D(n8288), .CK(CLK), .Q(net254140), .QN(
        n37011) );
  DFF_X1 \DRAM_mem_reg[30][12]  ( .D(n8287), .CK(CLK), .Q(net254139), .QN(
        n37010) );
  DFF_X1 \DRAM_mem_reg[30][11]  ( .D(n8286), .CK(CLK), .Q(net254138), .QN(
        n37009) );
  DFF_X1 \DRAM_mem_reg[30][10]  ( .D(n8285), .CK(CLK), .Q(net254137), .QN(
        n37008) );
  DFF_X1 \DRAM_mem_reg[30][9]  ( .D(n8284), .CK(CLK), .Q(net254136), .QN(
        n37007) );
  DFF_X1 \DRAM_mem_reg[30][8]  ( .D(n8283), .CK(CLK), .Q(net254135), .QN(
        n37006) );
  DFF_X1 \DRAM_mem_reg[30][7]  ( .D(n8282), .CK(CLK), .Q(net254134), .QN(
        n37005) );
  DFF_X1 \DRAM_mem_reg[30][6]  ( .D(n8281), .CK(CLK), .Q(net254133), .QN(
        n37004) );
  DFF_X1 \DRAM_mem_reg[30][5]  ( .D(n8280), .CK(CLK), .Q(net254132), .QN(
        n37003) );
  DFF_X1 \DRAM_mem_reg[30][4]  ( .D(n8279), .CK(CLK), .Q(net254131), .QN(
        n37002) );
  DFF_X1 \DRAM_mem_reg[30][3]  ( .D(n8278), .CK(CLK), .Q(net254130), .QN(
        n37001) );
  DFF_X1 \DRAM_mem_reg[30][2]  ( .D(n8277), .CK(CLK), .Q(net254129), .QN(
        n37000) );
  DFF_X1 \DRAM_mem_reg[30][1]  ( .D(n8276), .CK(CLK), .Q(net254128), .QN(
        n36999) );
  DFF_X1 \DRAM_mem_reg[30][0]  ( .D(n8275), .CK(CLK), .Q(net254127), .QN(
        n36998) );
  DFF_X1 \DRAM_mem_reg[31][31]  ( .D(n8274), .CK(CLK), .QN(n35408) );
  DFF_X1 \DRAM_mem_reg[31][30]  ( .D(n8273), .CK(CLK), .QN(n35399) );
  DFF_X1 \DRAM_mem_reg[31][29]  ( .D(n8272), .CK(CLK), .QN(n35390) );
  DFF_X1 \DRAM_mem_reg[31][28]  ( .D(n8271), .CK(CLK), .QN(n35381) );
  DFF_X1 \DRAM_mem_reg[31][27]  ( .D(n8270), .CK(CLK), .QN(n35372) );
  DFF_X1 \DRAM_mem_reg[31][26]  ( .D(n8269), .CK(CLK), .QN(n35363) );
  DFF_X1 \DRAM_mem_reg[31][25]  ( .D(n8268), .CK(CLK), .QN(n35354) );
  DFF_X1 \DRAM_mem_reg[31][24]  ( .D(n8267), .CK(CLK), .QN(n35345) );
  DFF_X1 \DRAM_mem_reg[31][23]  ( .D(n8266), .CK(CLK), .QN(n35612) );
  DFF_X1 \DRAM_mem_reg[31][22]  ( .D(n8265), .CK(CLK), .QN(n35610) );
  DFF_X1 \DRAM_mem_reg[31][21]  ( .D(n8264), .CK(CLK), .QN(n35608) );
  DFF_X1 \DRAM_mem_reg[31][20]  ( .D(n8263), .CK(CLK), .QN(n35606) );
  DFF_X1 \DRAM_mem_reg[31][19]  ( .D(n8262), .CK(CLK), .QN(n35604) );
  DFF_X1 \DRAM_mem_reg[31][18]  ( .D(n8261), .CK(CLK), .QN(n35602) );
  DFF_X1 \DRAM_mem_reg[31][17]  ( .D(n8260), .CK(CLK), .QN(n35600) );
  DFF_X1 \DRAM_mem_reg[31][16]  ( .D(n8259), .CK(CLK), .QN(n35598) );
  DFF_X1 \DRAM_mem_reg[31][15]  ( .D(n8258), .CK(CLK), .QN(n35596) );
  DFF_X1 \DRAM_mem_reg[31][14]  ( .D(n8257), .CK(CLK), .QN(n35594) );
  DFF_X1 \DRAM_mem_reg[31][13]  ( .D(n8256), .CK(CLK), .QN(n35592) );
  DFF_X1 \DRAM_mem_reg[31][12]  ( .D(n8255), .CK(CLK), .QN(n35590) );
  DFF_X1 \DRAM_mem_reg[31][11]  ( .D(n8254), .CK(CLK), .QN(n35588) );
  DFF_X1 \DRAM_mem_reg[31][10]  ( .D(n8253), .CK(CLK), .QN(n35586) );
  DFF_X1 \DRAM_mem_reg[31][9]  ( .D(n8252), .CK(CLK), .QN(n35584) );
  DFF_X1 \DRAM_mem_reg[31][8]  ( .D(n8251), .CK(CLK), .QN(n35582) );
  DFF_X1 \DRAM_mem_reg[31][7]  ( .D(n8250), .CK(CLK), .QN(n35580) );
  DFF_X1 \DRAM_mem_reg[31][6]  ( .D(n8249), .CK(CLK), .QN(n35578) );
  DFF_X1 \DRAM_mem_reg[31][5]  ( .D(n8248), .CK(CLK), .QN(n35576) );
  DFF_X1 \DRAM_mem_reg[31][4]  ( .D(n8247), .CK(CLK), .QN(n35574) );
  DFF_X1 \DRAM_mem_reg[31][3]  ( .D(n8246), .CK(CLK), .QN(n35572) );
  DFF_X1 \DRAM_mem_reg[31][2]  ( .D(n8245), .CK(CLK), .QN(n35570) );
  DFF_X1 \DRAM_mem_reg[31][1]  ( .D(n8244), .CK(CLK), .QN(n35568) );
  DFF_X1 \DRAM_mem_reg[31][0]  ( .D(n8243), .CK(CLK), .QN(n35566) );
  DFF_X1 \DRAM_mem_reg[32][31]  ( .D(n8242), .CK(CLK), .QN(n36205) );
  DFF_X1 \DRAM_mem_reg[32][30]  ( .D(n8241), .CK(CLK), .QN(n36204) );
  DFF_X1 \DRAM_mem_reg[32][29]  ( .D(n8240), .CK(CLK), .QN(n36203) );
  DFF_X1 \DRAM_mem_reg[32][28]  ( .D(n8239), .CK(CLK), .QN(n36202) );
  DFF_X1 \DRAM_mem_reg[32][27]  ( .D(n8238), .CK(CLK), .QN(n36201) );
  DFF_X1 \DRAM_mem_reg[32][26]  ( .D(n8237), .CK(CLK), .QN(n36200) );
  DFF_X1 \DRAM_mem_reg[32][25]  ( .D(n8236), .CK(CLK), .QN(n36199) );
  DFF_X1 \DRAM_mem_reg[32][24]  ( .D(n8235), .CK(CLK), .QN(n36198) );
  DFF_X1 \DRAM_mem_reg[32][23]  ( .D(n8234), .CK(CLK), .QN(n36317) );
  DFF_X1 \DRAM_mem_reg[32][22]  ( .D(n8233), .CK(CLK), .QN(n36316) );
  DFF_X1 \DRAM_mem_reg[32][21]  ( .D(n8232), .CK(CLK), .QN(n36315) );
  DFF_X1 \DRAM_mem_reg[32][20]  ( .D(n8231), .CK(CLK), .QN(n36314) );
  DFF_X1 \DRAM_mem_reg[32][19]  ( .D(n8230), .CK(CLK), .QN(n36313) );
  DFF_X1 \DRAM_mem_reg[32][18]  ( .D(n8229), .CK(CLK), .QN(n36312) );
  DFF_X1 \DRAM_mem_reg[32][17]  ( .D(n8228), .CK(CLK), .QN(n36311) );
  DFF_X1 \DRAM_mem_reg[32][16]  ( .D(n8227), .CK(CLK), .QN(n36310) );
  DFF_X1 \DRAM_mem_reg[32][15]  ( .D(n8226), .CK(CLK), .QN(n36309) );
  DFF_X1 \DRAM_mem_reg[32][14]  ( .D(n8225), .CK(CLK), .QN(n36308) );
  DFF_X1 \DRAM_mem_reg[32][13]  ( .D(n8224), .CK(CLK), .QN(n36307) );
  DFF_X1 \DRAM_mem_reg[32][12]  ( .D(n8223), .CK(CLK), .QN(n36306) );
  DFF_X1 \DRAM_mem_reg[32][11]  ( .D(n8222), .CK(CLK), .QN(n36305) );
  DFF_X1 \DRAM_mem_reg[32][10]  ( .D(n8221), .CK(CLK), .QN(n36304) );
  DFF_X1 \DRAM_mem_reg[32][9]  ( .D(n8220), .CK(CLK), .QN(n36303) );
  DFF_X1 \DRAM_mem_reg[32][8]  ( .D(n8219), .CK(CLK), .QN(n36302) );
  DFF_X1 \DRAM_mem_reg[32][7]  ( .D(n8218), .CK(CLK), .QN(n36301) );
  DFF_X1 \DRAM_mem_reg[32][6]  ( .D(n8217), .CK(CLK), .QN(n36300) );
  DFF_X1 \DRAM_mem_reg[32][5]  ( .D(n8216), .CK(CLK), .QN(n36299) );
  DFF_X1 \DRAM_mem_reg[32][4]  ( .D(n8215), .CK(CLK), .QN(n36298) );
  DFF_X1 \DRAM_mem_reg[32][3]  ( .D(n8214), .CK(CLK), .QN(n36297) );
  DFF_X1 \DRAM_mem_reg[32][2]  ( .D(n8213), .CK(CLK), .QN(n36296) );
  DFF_X1 \DRAM_mem_reg[32][1]  ( .D(n8212), .CK(CLK), .QN(n36295) );
  DFF_X1 \DRAM_mem_reg[32][0]  ( .D(n8211), .CK(CLK), .QN(n36294) );
  DFF_X1 \DRAM_mem_reg[33][31]  ( .D(n8210), .CK(CLK), .Q(net254126), .QN(
        n36757) );
  DFF_X1 \DRAM_mem_reg[33][30]  ( .D(n8209), .CK(CLK), .Q(net254125), .QN(
        n36756) );
  DFF_X1 \DRAM_mem_reg[33][29]  ( .D(n8208), .CK(CLK), .Q(net254124), .QN(
        n36755) );
  DFF_X1 \DRAM_mem_reg[33][28]  ( .D(n8207), .CK(CLK), .Q(net254123), .QN(
        n36754) );
  DFF_X1 \DRAM_mem_reg[33][27]  ( .D(n8206), .CK(CLK), .Q(net254122), .QN(
        n36753) );
  DFF_X1 \DRAM_mem_reg[33][26]  ( .D(n8205), .CK(CLK), .Q(net254121), .QN(
        n36752) );
  DFF_X1 \DRAM_mem_reg[33][25]  ( .D(n8204), .CK(CLK), .Q(net254120), .QN(
        n36751) );
  DFF_X1 \DRAM_mem_reg[33][24]  ( .D(n8203), .CK(CLK), .Q(net254119), .QN(
        n36750) );
  DFF_X1 \DRAM_mem_reg[33][23]  ( .D(n8202), .CK(CLK), .Q(net254118), .QN(
        n36997) );
  DFF_X1 \DRAM_mem_reg[33][22]  ( .D(n8201), .CK(CLK), .Q(net254117), .QN(
        n36996) );
  DFF_X1 \DRAM_mem_reg[33][21]  ( .D(n8200), .CK(CLK), .Q(net254116), .QN(
        n36995) );
  DFF_X1 \DRAM_mem_reg[33][20]  ( .D(n8199), .CK(CLK), .Q(net254115), .QN(
        n36994) );
  DFF_X1 \DRAM_mem_reg[33][19]  ( .D(n8198), .CK(CLK), .Q(net254114), .QN(
        n36993) );
  DFF_X1 \DRAM_mem_reg[33][18]  ( .D(n8197), .CK(CLK), .Q(net254113), .QN(
        n36992) );
  DFF_X1 \DRAM_mem_reg[33][17]  ( .D(n8196), .CK(CLK), .Q(net254112), .QN(
        n36991) );
  DFF_X1 \DRAM_mem_reg[33][16]  ( .D(n8195), .CK(CLK), .Q(net254111), .QN(
        n36990) );
  DFF_X1 \DRAM_mem_reg[33][15]  ( .D(n8194), .CK(CLK), .Q(net254110), .QN(
        n36989) );
  DFF_X1 \DRAM_mem_reg[33][14]  ( .D(n8193), .CK(CLK), .Q(net254109), .QN(
        n36988) );
  DFF_X1 \DRAM_mem_reg[33][13]  ( .D(n8192), .CK(CLK), .Q(net254108), .QN(
        n36987) );
  DFF_X1 \DRAM_mem_reg[33][12]  ( .D(n8191), .CK(CLK), .Q(net254107), .QN(
        n36986) );
  DFF_X1 \DRAM_mem_reg[33][11]  ( .D(n8190), .CK(CLK), .Q(net254106), .QN(
        n36985) );
  DFF_X1 \DRAM_mem_reg[33][10]  ( .D(n8189), .CK(CLK), .Q(net254105), .QN(
        n36984) );
  DFF_X1 \DRAM_mem_reg[33][9]  ( .D(n8188), .CK(CLK), .Q(net254104), .QN(
        n36983) );
  DFF_X1 \DRAM_mem_reg[33][8]  ( .D(n8187), .CK(CLK), .Q(net254103), .QN(
        n36982) );
  DFF_X1 \DRAM_mem_reg[33][7]  ( .D(n8186), .CK(CLK), .Q(net254102), .QN(
        n36981) );
  DFF_X1 \DRAM_mem_reg[33][6]  ( .D(n8185), .CK(CLK), .Q(net254101), .QN(
        n36980) );
  DFF_X1 \DRAM_mem_reg[33][5]  ( .D(n8184), .CK(CLK), .Q(net254100), .QN(
        n36979) );
  DFF_X1 \DRAM_mem_reg[33][4]  ( .D(n8183), .CK(CLK), .Q(net254099), .QN(
        n36978) );
  DFF_X1 \DRAM_mem_reg[33][3]  ( .D(n8182), .CK(CLK), .Q(net254098), .QN(
        n36977) );
  DFF_X1 \DRAM_mem_reg[33][2]  ( .D(n8181), .CK(CLK), .Q(net254097), .QN(
        n36976) );
  DFF_X1 \DRAM_mem_reg[33][1]  ( .D(n8180), .CK(CLK), .Q(net254096), .QN(
        n36975) );
  DFF_X1 \DRAM_mem_reg[33][0]  ( .D(n8179), .CK(CLK), .Q(net254095), .QN(
        n36974) );
  DFF_X1 \DRAM_mem_reg[34][31]  ( .D(n8178), .CK(CLK), .QN(n35173) );
  DFF_X1 \DRAM_mem_reg[34][30]  ( .D(n8177), .CK(CLK), .QN(n35172) );
  DFF_X1 \DRAM_mem_reg[34][29]  ( .D(n8176), .CK(CLK), .QN(n35171) );
  DFF_X1 \DRAM_mem_reg[34][28]  ( .D(n8175), .CK(CLK), .QN(n35170) );
  DFF_X1 \DRAM_mem_reg[34][27]  ( .D(n8174), .CK(CLK), .QN(n35169) );
  DFF_X1 \DRAM_mem_reg[34][26]  ( .D(n8173), .CK(CLK), .QN(n35168) );
  DFF_X1 \DRAM_mem_reg[34][25]  ( .D(n8172), .CK(CLK), .QN(n35167) );
  DFF_X1 \DRAM_mem_reg[34][24]  ( .D(n8171), .CK(CLK), .QN(n35166) );
  DFF_X1 \DRAM_mem_reg[34][23]  ( .D(n8170), .CK(CLK), .QN(n35269) );
  DFF_X1 \DRAM_mem_reg[34][22]  ( .D(n8169), .CK(CLK), .QN(n35268) );
  DFF_X1 \DRAM_mem_reg[34][21]  ( .D(n8168), .CK(CLK), .QN(n35267) );
  DFF_X1 \DRAM_mem_reg[34][20]  ( .D(n8167), .CK(CLK), .QN(n35266) );
  DFF_X1 \DRAM_mem_reg[34][19]  ( .D(n8166), .CK(CLK), .QN(n35265) );
  DFF_X1 \DRAM_mem_reg[34][18]  ( .D(n8165), .CK(CLK), .QN(n35264) );
  DFF_X1 \DRAM_mem_reg[34][17]  ( .D(n8164), .CK(CLK), .QN(n35263) );
  DFF_X1 \DRAM_mem_reg[34][16]  ( .D(n8163), .CK(CLK), .QN(n35262) );
  DFF_X1 \DRAM_mem_reg[34][15]  ( .D(n8162), .CK(CLK), .QN(n35261) );
  DFF_X1 \DRAM_mem_reg[34][14]  ( .D(n8161), .CK(CLK), .QN(n35260) );
  DFF_X1 \DRAM_mem_reg[34][13]  ( .D(n8160), .CK(CLK), .QN(n35259) );
  DFF_X1 \DRAM_mem_reg[34][12]  ( .D(n8159), .CK(CLK), .QN(n35258) );
  DFF_X1 \DRAM_mem_reg[34][11]  ( .D(n8158), .CK(CLK), .QN(n35257) );
  DFF_X1 \DRAM_mem_reg[34][10]  ( .D(n8157), .CK(CLK), .QN(n35256) );
  DFF_X1 \DRAM_mem_reg[34][9]  ( .D(n8156), .CK(CLK), .QN(n35255) );
  DFF_X1 \DRAM_mem_reg[34][8]  ( .D(n8155), .CK(CLK), .QN(n35254) );
  DFF_X1 \DRAM_mem_reg[34][7]  ( .D(n8154), .CK(CLK), .QN(n35253) );
  DFF_X1 \DRAM_mem_reg[34][6]  ( .D(n8153), .CK(CLK), .QN(n35252) );
  DFF_X1 \DRAM_mem_reg[34][5]  ( .D(n8152), .CK(CLK), .QN(n35251) );
  DFF_X1 \DRAM_mem_reg[34][4]  ( .D(n8151), .CK(CLK), .QN(n35250) );
  DFF_X1 \DRAM_mem_reg[34][3]  ( .D(n8150), .CK(CLK), .QN(n35249) );
  DFF_X1 \DRAM_mem_reg[34][2]  ( .D(n8149), .CK(CLK), .QN(n35248) );
  DFF_X1 \DRAM_mem_reg[34][1]  ( .D(n8148), .CK(CLK), .QN(n35247) );
  DFF_X1 \DRAM_mem_reg[34][0]  ( .D(n8147), .CK(CLK), .QN(n35246) );
  DFF_X1 \DRAM_mem_reg[35][31]  ( .D(n8146), .CK(CLK), .QN(n35923) );
  DFF_X1 \DRAM_mem_reg[35][30]  ( .D(n8145), .CK(CLK), .QN(n35914) );
  DFF_X1 \DRAM_mem_reg[35][29]  ( .D(n8144), .CK(CLK), .QN(n35905) );
  DFF_X1 \DRAM_mem_reg[35][28]  ( .D(n8143), .CK(CLK), .QN(n35896) );
  DFF_X1 \DRAM_mem_reg[35][27]  ( .D(n8142), .CK(CLK), .QN(n35887) );
  DFF_X1 \DRAM_mem_reg[35][26]  ( .D(n8141), .CK(CLK), .QN(n35878) );
  DFF_X1 \DRAM_mem_reg[35][25]  ( .D(n8140), .CK(CLK), .QN(n35869) );
  DFF_X1 \DRAM_mem_reg[35][24]  ( .D(n8139), .CK(CLK), .QN(n35860) );
  DFF_X1 \DRAM_mem_reg[35][23]  ( .D(n8138), .CK(CLK), .QN(n36077) );
  DFF_X1 \DRAM_mem_reg[35][22]  ( .D(n8137), .CK(CLK), .QN(n36075) );
  DFF_X1 \DRAM_mem_reg[35][21]  ( .D(n8136), .CK(CLK), .QN(n36073) );
  DFF_X1 \DRAM_mem_reg[35][20]  ( .D(n8135), .CK(CLK), .QN(n36071) );
  DFF_X1 \DRAM_mem_reg[35][19]  ( .D(n8134), .CK(CLK), .QN(n36069) );
  DFF_X1 \DRAM_mem_reg[35][18]  ( .D(n8133), .CK(CLK), .QN(n36067) );
  DFF_X1 \DRAM_mem_reg[35][17]  ( .D(n8132), .CK(CLK), .QN(n36065) );
  DFF_X1 \DRAM_mem_reg[35][16]  ( .D(n8131), .CK(CLK), .QN(n36063) );
  DFF_X1 \DRAM_mem_reg[35][15]  ( .D(n8130), .CK(CLK), .QN(n36061) );
  DFF_X1 \DRAM_mem_reg[35][14]  ( .D(n8129), .CK(CLK), .QN(n36059) );
  DFF_X1 \DRAM_mem_reg[35][13]  ( .D(n8128), .CK(CLK), .QN(n36057) );
  DFF_X1 \DRAM_mem_reg[35][12]  ( .D(n8127), .CK(CLK), .QN(n36055) );
  DFF_X1 \DRAM_mem_reg[35][11]  ( .D(n8126), .CK(CLK), .QN(n36053) );
  DFF_X1 \DRAM_mem_reg[35][10]  ( .D(n8125), .CK(CLK), .QN(n36051) );
  DFF_X1 \DRAM_mem_reg[35][9]  ( .D(n8124), .CK(CLK), .QN(n36049) );
  DFF_X1 \DRAM_mem_reg[35][8]  ( .D(n8123), .CK(CLK), .QN(n36047) );
  DFF_X1 \DRAM_mem_reg[35][7]  ( .D(n8122), .CK(CLK), .QN(n36045) );
  DFF_X1 \DRAM_mem_reg[35][6]  ( .D(n8121), .CK(CLK), .QN(n36043) );
  DFF_X1 \DRAM_mem_reg[35][5]  ( .D(n8120), .CK(CLK), .QN(n36041) );
  DFF_X1 \DRAM_mem_reg[35][4]  ( .D(n8119), .CK(CLK), .QN(n36039) );
  DFF_X1 \DRAM_mem_reg[35][3]  ( .D(n8118), .CK(CLK), .QN(n36037) );
  DFF_X1 \DRAM_mem_reg[35][2]  ( .D(n8117), .CK(CLK), .QN(n36035) );
  DFF_X1 \DRAM_mem_reg[35][1]  ( .D(n8116), .CK(CLK), .QN(n36033) );
  DFF_X1 \DRAM_mem_reg[35][0]  ( .D(n8115), .CK(CLK), .QN(n36031) );
  DFF_X1 \DRAM_mem_reg[36][31]  ( .D(n8114), .CK(CLK), .Q(net254094), .QN(
        n37141) );
  DFF_X1 \DRAM_mem_reg[36][30]  ( .D(n8113), .CK(CLK), .Q(net254093), .QN(
        n37140) );
  DFF_X1 \DRAM_mem_reg[36][29]  ( .D(n8112), .CK(CLK), .Q(net254092), .QN(
        n37139) );
  DFF_X1 \DRAM_mem_reg[36][28]  ( .D(n8111), .CK(CLK), .Q(net254091), .QN(
        n37138) );
  DFF_X1 \DRAM_mem_reg[36][27]  ( .D(n8110), .CK(CLK), .Q(net254090), .QN(
        n37137) );
  DFF_X1 \DRAM_mem_reg[36][26]  ( .D(n8109), .CK(CLK), .Q(net254089), .QN(
        n37136) );
  DFF_X1 \DRAM_mem_reg[36][25]  ( .D(n8108), .CK(CLK), .Q(net254088), .QN(
        n37135) );
  DFF_X1 \DRAM_mem_reg[36][24]  ( .D(n8107), .CK(CLK), .Q(net254087), .QN(
        n37134) );
  DFF_X1 \DRAM_mem_reg[36][23]  ( .D(n8106), .CK(CLK), .Q(net254086), .QN(
        n37381) );
  DFF_X1 \DRAM_mem_reg[36][22]  ( .D(n8105), .CK(CLK), .Q(net254085), .QN(
        n37380) );
  DFF_X1 \DRAM_mem_reg[36][21]  ( .D(n8104), .CK(CLK), .Q(net254084), .QN(
        n37379) );
  DFF_X1 \DRAM_mem_reg[36][20]  ( .D(n8103), .CK(CLK), .Q(net254083), .QN(
        n37378) );
  DFF_X1 \DRAM_mem_reg[36][19]  ( .D(n8102), .CK(CLK), .Q(net254082), .QN(
        n37377) );
  DFF_X1 \DRAM_mem_reg[36][18]  ( .D(n8101), .CK(CLK), .Q(net254081), .QN(
        n37376) );
  DFF_X1 \DRAM_mem_reg[36][17]  ( .D(n8100), .CK(CLK), .Q(net254080), .QN(
        n37375) );
  DFF_X1 \DRAM_mem_reg[36][16]  ( .D(n8099), .CK(CLK), .Q(net254079), .QN(
        n37374) );
  DFF_X1 \DRAM_mem_reg[36][15]  ( .D(n8098), .CK(CLK), .Q(net254078), .QN(
        n37373) );
  DFF_X1 \DRAM_mem_reg[36][14]  ( .D(n8097), .CK(CLK), .Q(net254077), .QN(
        n37372) );
  DFF_X1 \DRAM_mem_reg[36][13]  ( .D(n8096), .CK(CLK), .Q(net254076), .QN(
        n37371) );
  DFF_X1 \DRAM_mem_reg[36][12]  ( .D(n8095), .CK(CLK), .Q(net254075), .QN(
        n37370) );
  DFF_X1 \DRAM_mem_reg[36][11]  ( .D(n8094), .CK(CLK), .Q(net254074), .QN(
        n37369) );
  DFF_X1 \DRAM_mem_reg[36][10]  ( .D(n8093), .CK(CLK), .Q(net254073), .QN(
        n37368) );
  DFF_X1 \DRAM_mem_reg[36][9]  ( .D(n8092), .CK(CLK), .Q(net254072), .QN(
        n37367) );
  DFF_X1 \DRAM_mem_reg[36][8]  ( .D(n8091), .CK(CLK), .Q(net254071), .QN(
        n37366) );
  DFF_X1 \DRAM_mem_reg[36][7]  ( .D(n8090), .CK(CLK), .Q(net254070), .QN(
        n37365) );
  DFF_X1 \DRAM_mem_reg[36][6]  ( .D(n8089), .CK(CLK), .Q(net254069), .QN(
        n37364) );
  DFF_X1 \DRAM_mem_reg[36][5]  ( .D(n8088), .CK(CLK), .Q(net254068), .QN(
        n37363) );
  DFF_X1 \DRAM_mem_reg[36][4]  ( .D(n8087), .CK(CLK), .Q(net254067), .QN(
        n37362) );
  DFF_X1 \DRAM_mem_reg[36][3]  ( .D(n8086), .CK(CLK), .Q(net254066), .QN(
        n37361) );
  DFF_X1 \DRAM_mem_reg[36][2]  ( .D(n8085), .CK(CLK), .Q(net254065), .QN(
        n37360) );
  DFF_X1 \DRAM_mem_reg[36][1]  ( .D(n8084), .CK(CLK), .Q(net254064), .QN(
        n37359) );
  DFF_X1 \DRAM_mem_reg[36][0]  ( .D(n8083), .CK(CLK), .Q(net254063), .QN(
        n37358) );
  DFF_X1 \DRAM_mem_reg[37][31]  ( .D(n8082), .CK(CLK), .QN(n36434) );
  DFF_X1 \DRAM_mem_reg[37][30]  ( .D(n8081), .CK(CLK), .QN(n36425) );
  DFF_X1 \DRAM_mem_reg[37][29]  ( .D(n8080), .CK(CLK), .QN(n36416) );
  DFF_X1 \DRAM_mem_reg[37][28]  ( .D(n8079), .CK(CLK), .QN(n36407) );
  DFF_X1 \DRAM_mem_reg[37][27]  ( .D(n8078), .CK(CLK), .QN(n36398) );
  DFF_X1 \DRAM_mem_reg[37][26]  ( .D(n8077), .CK(CLK), .QN(n36389) );
  DFF_X1 \DRAM_mem_reg[37][25]  ( .D(n8076), .CK(CLK), .QN(n36380) );
  DFF_X1 \DRAM_mem_reg[37][24]  ( .D(n8075), .CK(CLK), .QN(n36371) );
  DFF_X1 \DRAM_mem_reg[37][23]  ( .D(n8074), .CK(CLK), .QN(n36533) );
  DFF_X1 \DRAM_mem_reg[37][22]  ( .D(n8073), .CK(CLK), .QN(n36529) );
  DFF_X1 \DRAM_mem_reg[37][21]  ( .D(n8072), .CK(CLK), .QN(n36525) );
  DFF_X1 \DRAM_mem_reg[37][20]  ( .D(n8071), .CK(CLK), .QN(n36521) );
  DFF_X1 \DRAM_mem_reg[37][19]  ( .D(n8070), .CK(CLK), .QN(n36517) );
  DFF_X1 \DRAM_mem_reg[37][18]  ( .D(n8069), .CK(CLK), .QN(n36513) );
  DFF_X1 \DRAM_mem_reg[37][17]  ( .D(n8068), .CK(CLK), .QN(n36509) );
  DFF_X1 \DRAM_mem_reg[37][16]  ( .D(n8067), .CK(CLK), .QN(n36505) );
  DFF_X1 \DRAM_mem_reg[37][15]  ( .D(n8066), .CK(CLK), .QN(n36501) );
  DFF_X1 \DRAM_mem_reg[37][14]  ( .D(n8065), .CK(CLK), .QN(n36497) );
  DFF_X1 \DRAM_mem_reg[37][13]  ( .D(n8064), .CK(CLK), .QN(n36493) );
  DFF_X1 \DRAM_mem_reg[37][12]  ( .D(n8063), .CK(CLK), .QN(n36489) );
  DFF_X1 \DRAM_mem_reg[37][11]  ( .D(n8062), .CK(CLK), .QN(n36485) );
  DFF_X1 \DRAM_mem_reg[37][10]  ( .D(n8061), .CK(CLK), .QN(n36481) );
  DFF_X1 \DRAM_mem_reg[37][9]  ( .D(n8060), .CK(CLK), .QN(n36477) );
  DFF_X1 \DRAM_mem_reg[37][8]  ( .D(n8059), .CK(CLK), .QN(n36473) );
  DFF_X1 \DRAM_mem_reg[37][7]  ( .D(n8058), .CK(CLK), .QN(n36469) );
  DFF_X1 \DRAM_mem_reg[37][6]  ( .D(n8057), .CK(CLK), .QN(n36465) );
  DFF_X1 \DRAM_mem_reg[37][5]  ( .D(n8056), .CK(CLK), .QN(n36461) );
  DFF_X1 \DRAM_mem_reg[37][4]  ( .D(n8055), .CK(CLK), .QN(n36457) );
  DFF_X1 \DRAM_mem_reg[37][3]  ( .D(n8054), .CK(CLK), .QN(n36453) );
  DFF_X1 \DRAM_mem_reg[37][2]  ( .D(n8053), .CK(CLK), .QN(n36449) );
  DFF_X1 \DRAM_mem_reg[37][1]  ( .D(n8052), .CK(CLK), .QN(n36445) );
  DFF_X1 \DRAM_mem_reg[37][0]  ( .D(n8051), .CK(CLK), .QN(n36441) );
  DFF_X1 \DRAM_mem_reg[38][31]  ( .D(n8050), .CK(CLK), .Q(net254062), .QN(
        n36749) );
  DFF_X1 \DRAM_mem_reg[38][30]  ( .D(n8049), .CK(CLK), .Q(net254061), .QN(
        n36748) );
  DFF_X1 \DRAM_mem_reg[38][29]  ( .D(n8048), .CK(CLK), .Q(net254060), .QN(
        n36747) );
  DFF_X1 \DRAM_mem_reg[38][28]  ( .D(n8047), .CK(CLK), .Q(net254059), .QN(
        n36746) );
  DFF_X1 \DRAM_mem_reg[38][27]  ( .D(n8046), .CK(CLK), .Q(net254058), .QN(
        n36745) );
  DFF_X1 \DRAM_mem_reg[38][26]  ( .D(n8045), .CK(CLK), .Q(net254057), .QN(
        n36744) );
  DFF_X1 \DRAM_mem_reg[38][25]  ( .D(n8044), .CK(CLK), .Q(net254056), .QN(
        n36743) );
  DFF_X1 \DRAM_mem_reg[38][24]  ( .D(n8043), .CK(CLK), .Q(net254055), .QN(
        n36742) );
  DFF_X1 \DRAM_mem_reg[38][23]  ( .D(n8042), .CK(CLK), .Q(net254054), .QN(
        n36973) );
  DFF_X1 \DRAM_mem_reg[38][22]  ( .D(n8041), .CK(CLK), .Q(net254053), .QN(
        n36972) );
  DFF_X1 \DRAM_mem_reg[38][21]  ( .D(n8040), .CK(CLK), .Q(net254052), .QN(
        n36971) );
  DFF_X1 \DRAM_mem_reg[38][20]  ( .D(n8039), .CK(CLK), .Q(net254051), .QN(
        n36970) );
  DFF_X1 \DRAM_mem_reg[38][19]  ( .D(n8038), .CK(CLK), .Q(net254050), .QN(
        n36969) );
  DFF_X1 \DRAM_mem_reg[38][18]  ( .D(n8037), .CK(CLK), .Q(net254049), .QN(
        n36968) );
  DFF_X1 \DRAM_mem_reg[38][17]  ( .D(n8036), .CK(CLK), .Q(net254048), .QN(
        n36967) );
  DFF_X1 \DRAM_mem_reg[38][16]  ( .D(n8035), .CK(CLK), .Q(net254047), .QN(
        n36966) );
  DFF_X1 \DRAM_mem_reg[38][15]  ( .D(n8034), .CK(CLK), .Q(net254046), .QN(
        n36965) );
  DFF_X1 \DRAM_mem_reg[38][14]  ( .D(n8033), .CK(CLK), .Q(net254045), .QN(
        n36964) );
  DFF_X1 \DRAM_mem_reg[38][13]  ( .D(n8032), .CK(CLK), .Q(net254044), .QN(
        n36963) );
  DFF_X1 \DRAM_mem_reg[38][12]  ( .D(n8031), .CK(CLK), .Q(net254043), .QN(
        n36962) );
  DFF_X1 \DRAM_mem_reg[38][11]  ( .D(n8030), .CK(CLK), .Q(net254042), .QN(
        n36961) );
  DFF_X1 \DRAM_mem_reg[38][10]  ( .D(n8029), .CK(CLK), .Q(net254041), .QN(
        n36960) );
  DFF_X1 \DRAM_mem_reg[38][9]  ( .D(n8028), .CK(CLK), .Q(net254040), .QN(
        n36959) );
  DFF_X1 \DRAM_mem_reg[38][8]  ( .D(n8027), .CK(CLK), .Q(net254039), .QN(
        n36958) );
  DFF_X1 \DRAM_mem_reg[38][7]  ( .D(n8026), .CK(CLK), .Q(net254038), .QN(
        n36957) );
  DFF_X1 \DRAM_mem_reg[38][6]  ( .D(n8025), .CK(CLK), .Q(net254037), .QN(
        n36956) );
  DFF_X1 \DRAM_mem_reg[38][5]  ( .D(n8024), .CK(CLK), .Q(net254036), .QN(
        n36955) );
  DFF_X1 \DRAM_mem_reg[38][4]  ( .D(n8023), .CK(CLK), .Q(net254035), .QN(
        n36954) );
  DFF_X1 \DRAM_mem_reg[38][3]  ( .D(n8022), .CK(CLK), .Q(net254034), .QN(
        n36953) );
  DFF_X1 \DRAM_mem_reg[38][2]  ( .D(n8021), .CK(CLK), .Q(net254033), .QN(
        n36952) );
  DFF_X1 \DRAM_mem_reg[38][1]  ( .D(n8020), .CK(CLK), .Q(net254032), .QN(
        n36951) );
  DFF_X1 \DRAM_mem_reg[38][0]  ( .D(n8019), .CK(CLK), .Q(net254031), .QN(
        n36950) );
  DFF_X1 \DRAM_mem_reg[39][31]  ( .D(n8018), .CK(CLK), .QN(n35413) );
  DFF_X1 \DRAM_mem_reg[39][30]  ( .D(n8017), .CK(CLK), .QN(n35404) );
  DFF_X1 \DRAM_mem_reg[39][29]  ( .D(n8016), .CK(CLK), .QN(n35395) );
  DFF_X1 \DRAM_mem_reg[39][28]  ( .D(n8015), .CK(CLK), .QN(n35386) );
  DFF_X1 \DRAM_mem_reg[39][27]  ( .D(n8014), .CK(CLK), .QN(n35377) );
  DFF_X1 \DRAM_mem_reg[39][26]  ( .D(n8013), .CK(CLK), .QN(n35368) );
  DFF_X1 \DRAM_mem_reg[39][25]  ( .D(n8012), .CK(CLK), .QN(n35359) );
  DFF_X1 \DRAM_mem_reg[39][24]  ( .D(n8011), .CK(CLK), .QN(n35350) );
  DFF_X1 \DRAM_mem_reg[39][23]  ( .D(n8010), .CK(CLK), .QN(n35661) );
  DFF_X1 \DRAM_mem_reg[39][22]  ( .D(n8009), .CK(CLK), .QN(n35659) );
  DFF_X1 \DRAM_mem_reg[39][21]  ( .D(n8008), .CK(CLK), .QN(n35657) );
  DFF_X1 \DRAM_mem_reg[39][20]  ( .D(n8007), .CK(CLK), .QN(n35655) );
  DFF_X1 \DRAM_mem_reg[39][19]  ( .D(n8006), .CK(CLK), .QN(n35653) );
  DFF_X1 \DRAM_mem_reg[39][18]  ( .D(n8005), .CK(CLK), .QN(n35651) );
  DFF_X1 \DRAM_mem_reg[39][17]  ( .D(n8004), .CK(CLK), .QN(n35649) );
  DFF_X1 \DRAM_mem_reg[39][16]  ( .D(n8003), .CK(CLK), .QN(n35647) );
  DFF_X1 \DRAM_mem_reg[39][15]  ( .D(n8002), .CK(CLK), .QN(n35645) );
  DFF_X1 \DRAM_mem_reg[39][14]  ( .D(n8001), .CK(CLK), .QN(n35643) );
  DFF_X1 \DRAM_mem_reg[39][13]  ( .D(n8000), .CK(CLK), .QN(n35641) );
  DFF_X1 \DRAM_mem_reg[39][12]  ( .D(n7999), .CK(CLK), .QN(n35639) );
  DFF_X1 \DRAM_mem_reg[39][11]  ( .D(n7998), .CK(CLK), .QN(n35637) );
  DFF_X1 \DRAM_mem_reg[39][10]  ( .D(n7997), .CK(CLK), .QN(n35635) );
  DFF_X1 \DRAM_mem_reg[39][9]  ( .D(n7996), .CK(CLK), .QN(n35633) );
  DFF_X1 \DRAM_mem_reg[39][8]  ( .D(n7995), .CK(CLK), .QN(n35631) );
  DFF_X1 \DRAM_mem_reg[39][7]  ( .D(n7994), .CK(CLK), .QN(n35629) );
  DFF_X1 \DRAM_mem_reg[39][6]  ( .D(n7993), .CK(CLK), .QN(n35627) );
  DFF_X1 \DRAM_mem_reg[39][5]  ( .D(n7992), .CK(CLK), .QN(n35625) );
  DFF_X1 \DRAM_mem_reg[39][4]  ( .D(n7991), .CK(CLK), .QN(n35623) );
  DFF_X1 \DRAM_mem_reg[39][3]  ( .D(n7990), .CK(CLK), .QN(n35621) );
  DFF_X1 \DRAM_mem_reg[39][2]  ( .D(n7989), .CK(CLK), .QN(n35619) );
  DFF_X1 \DRAM_mem_reg[39][1]  ( .D(n7988), .CK(CLK), .QN(n35617) );
  DFF_X1 \DRAM_mem_reg[39][0]  ( .D(n7987), .CK(CLK), .QN(n35615) );
  DFF_X1 \DRAM_mem_reg[40][31]  ( .D(n7986), .CK(CLK), .QN(n35924) );
  DFF_X1 \DRAM_mem_reg[40][30]  ( .D(n7985), .CK(CLK), .QN(n35915) );
  DFF_X1 \DRAM_mem_reg[40][29]  ( .D(n7984), .CK(CLK), .QN(n35906) );
  DFF_X1 \DRAM_mem_reg[40][28]  ( .D(n7983), .CK(CLK), .QN(n35897) );
  DFF_X1 \DRAM_mem_reg[40][27]  ( .D(n7982), .CK(CLK), .QN(n35888) );
  DFF_X1 \DRAM_mem_reg[40][26]  ( .D(n7981), .CK(CLK), .QN(n35879) );
  DFF_X1 \DRAM_mem_reg[40][25]  ( .D(n7980), .CK(CLK), .QN(n35870) );
  DFF_X1 \DRAM_mem_reg[40][24]  ( .D(n7979), .CK(CLK), .QN(n35861) );
  DFF_X1 \DRAM_mem_reg[40][23]  ( .D(n7978), .CK(CLK), .QN(n36125) );
  DFF_X1 \DRAM_mem_reg[40][22]  ( .D(n7977), .CK(CLK), .QN(n36123) );
  DFF_X1 \DRAM_mem_reg[40][21]  ( .D(n7976), .CK(CLK), .QN(n36121) );
  DFF_X1 \DRAM_mem_reg[40][20]  ( .D(n7975), .CK(CLK), .QN(n36119) );
  DFF_X1 \DRAM_mem_reg[40][19]  ( .D(n7974), .CK(CLK), .QN(n36117) );
  DFF_X1 \DRAM_mem_reg[40][18]  ( .D(n7973), .CK(CLK), .QN(n36115) );
  DFF_X1 \DRAM_mem_reg[40][17]  ( .D(n7972), .CK(CLK), .QN(n36113) );
  DFF_X1 \DRAM_mem_reg[40][16]  ( .D(n7971), .CK(CLK), .QN(n36111) );
  DFF_X1 \DRAM_mem_reg[40][15]  ( .D(n7970), .CK(CLK), .QN(n36109) );
  DFF_X1 \DRAM_mem_reg[40][14]  ( .D(n7969), .CK(CLK), .QN(n36107) );
  DFF_X1 \DRAM_mem_reg[40][13]  ( .D(n7968), .CK(CLK), .QN(n36105) );
  DFF_X1 \DRAM_mem_reg[40][12]  ( .D(n7967), .CK(CLK), .QN(n36103) );
  DFF_X1 \DRAM_mem_reg[40][11]  ( .D(n7966), .CK(CLK), .QN(n36101) );
  DFF_X1 \DRAM_mem_reg[40][10]  ( .D(n7965), .CK(CLK), .QN(n36099) );
  DFF_X1 \DRAM_mem_reg[40][9]  ( .D(n7964), .CK(CLK), .QN(n36097) );
  DFF_X1 \DRAM_mem_reg[40][8]  ( .D(n7963), .CK(CLK), .QN(n36095) );
  DFF_X1 \DRAM_mem_reg[40][7]  ( .D(n7962), .CK(CLK), .QN(n36093) );
  DFF_X1 \DRAM_mem_reg[40][6]  ( .D(n7961), .CK(CLK), .QN(n36091) );
  DFF_X1 \DRAM_mem_reg[40][5]  ( .D(n7960), .CK(CLK), .QN(n36089) );
  DFF_X1 \DRAM_mem_reg[40][4]  ( .D(n7959), .CK(CLK), .QN(n36087) );
  DFF_X1 \DRAM_mem_reg[40][3]  ( .D(n7958), .CK(CLK), .QN(n36085) );
  DFF_X1 \DRAM_mem_reg[40][2]  ( .D(n7957), .CK(CLK), .QN(n36083) );
  DFF_X1 \DRAM_mem_reg[40][1]  ( .D(n7956), .CK(CLK), .QN(n36081) );
  DFF_X1 \DRAM_mem_reg[40][0]  ( .D(n7955), .CK(CLK), .QN(n36079) );
  DFF_X1 \DRAM_mem_reg[41][31]  ( .D(n7954), .CK(CLK), .Q(net254030), .QN(
        n37133) );
  DFF_X1 \DRAM_mem_reg[41][30]  ( .D(n7953), .CK(CLK), .Q(net254029), .QN(
        n37132) );
  DFF_X1 \DRAM_mem_reg[41][29]  ( .D(n7952), .CK(CLK), .Q(net254028), .QN(
        n37131) );
  DFF_X1 \DRAM_mem_reg[41][28]  ( .D(n7951), .CK(CLK), .Q(net254027), .QN(
        n37130) );
  DFF_X1 \DRAM_mem_reg[41][27]  ( .D(n7950), .CK(CLK), .Q(net254026), .QN(
        n37129) );
  DFF_X1 \DRAM_mem_reg[41][26]  ( .D(n7949), .CK(CLK), .Q(net254025), .QN(
        n37128) );
  DFF_X1 \DRAM_mem_reg[41][25]  ( .D(n7948), .CK(CLK), .Q(net254024), .QN(
        n37127) );
  DFF_X1 \DRAM_mem_reg[41][24]  ( .D(n7947), .CK(CLK), .Q(net254023), .QN(
        n37126) );
  DFF_X1 \DRAM_mem_reg[41][23]  ( .D(n7946), .CK(CLK), .Q(net254022), .QN(
        n37357) );
  DFF_X1 \DRAM_mem_reg[41][22]  ( .D(n7945), .CK(CLK), .Q(net254021), .QN(
        n37356) );
  DFF_X1 \DRAM_mem_reg[41][21]  ( .D(n7944), .CK(CLK), .Q(net254020), .QN(
        n37355) );
  DFF_X1 \DRAM_mem_reg[41][20]  ( .D(n7943), .CK(CLK), .Q(net254019), .QN(
        n37354) );
  DFF_X1 \DRAM_mem_reg[41][19]  ( .D(n7942), .CK(CLK), .Q(net254018), .QN(
        n37353) );
  DFF_X1 \DRAM_mem_reg[41][18]  ( .D(n7941), .CK(CLK), .Q(net254017), .QN(
        n37352) );
  DFF_X1 \DRAM_mem_reg[41][17]  ( .D(n7940), .CK(CLK), .Q(net254016), .QN(
        n37351) );
  DFF_X1 \DRAM_mem_reg[41][16]  ( .D(n7939), .CK(CLK), .Q(net254015), .QN(
        n37350) );
  DFF_X1 \DRAM_mem_reg[41][15]  ( .D(n7938), .CK(CLK), .Q(net254014), .QN(
        n37349) );
  DFF_X1 \DRAM_mem_reg[41][14]  ( .D(n7937), .CK(CLK), .Q(net254013), .QN(
        n37348) );
  DFF_X1 \DRAM_mem_reg[41][13]  ( .D(n7936), .CK(CLK), .Q(net254012), .QN(
        n37347) );
  DFF_X1 \DRAM_mem_reg[41][12]  ( .D(n7935), .CK(CLK), .Q(net254011), .QN(
        n37346) );
  DFF_X1 \DRAM_mem_reg[41][11]  ( .D(n7934), .CK(CLK), .Q(net254010), .QN(
        n37345) );
  DFF_X1 \DRAM_mem_reg[41][10]  ( .D(n7933), .CK(CLK), .Q(net254009), .QN(
        n37344) );
  DFF_X1 \DRAM_mem_reg[41][9]  ( .D(n7932), .CK(CLK), .Q(net254008), .QN(
        n37343) );
  DFF_X1 \DRAM_mem_reg[41][8]  ( .D(n7931), .CK(CLK), .Q(net254007), .QN(
        n37342) );
  DFF_X1 \DRAM_mem_reg[41][7]  ( .D(n7930), .CK(CLK), .Q(net254006), .QN(
        n37341) );
  DFF_X1 \DRAM_mem_reg[41][6]  ( .D(n7929), .CK(CLK), .Q(net254005), .QN(
        n37340) );
  DFF_X1 \DRAM_mem_reg[41][5]  ( .D(n7928), .CK(CLK), .Q(net254004), .QN(
        n37339) );
  DFF_X1 \DRAM_mem_reg[41][4]  ( .D(n7927), .CK(CLK), .Q(net254003), .QN(
        n37338) );
  DFF_X1 \DRAM_mem_reg[41][3]  ( .D(n7926), .CK(CLK), .Q(net254002), .QN(
        n37337) );
  DFF_X1 \DRAM_mem_reg[41][2]  ( .D(n7925), .CK(CLK), .Q(net254001), .QN(
        n37336) );
  DFF_X1 \DRAM_mem_reg[41][1]  ( .D(n7924), .CK(CLK), .Q(net254000), .QN(
        n37335) );
  DFF_X1 \DRAM_mem_reg[41][0]  ( .D(n7923), .CK(CLK), .Q(net253999), .QN(
        n37334) );
  DFF_X1 \DRAM_mem_reg[42][31]  ( .D(n7922), .CK(CLK), .QN(n36431) );
  DFF_X1 \DRAM_mem_reg[42][30]  ( .D(n7921), .CK(CLK), .QN(n36422) );
  DFF_X1 \DRAM_mem_reg[42][29]  ( .D(n7920), .CK(CLK), .QN(n36413) );
  DFF_X1 \DRAM_mem_reg[42][28]  ( .D(n7919), .CK(CLK), .QN(n36404) );
  DFF_X1 \DRAM_mem_reg[42][27]  ( .D(n7918), .CK(CLK), .QN(n36395) );
  DFF_X1 \DRAM_mem_reg[42][26]  ( .D(n7917), .CK(CLK), .QN(n36386) );
  DFF_X1 \DRAM_mem_reg[42][25]  ( .D(n7916), .CK(CLK), .QN(n36377) );
  DFF_X1 \DRAM_mem_reg[42][24]  ( .D(n7915), .CK(CLK), .QN(n36368) );
  DFF_X1 \DRAM_mem_reg[42][23]  ( .D(n7914), .CK(CLK), .QN(n36588) );
  DFF_X1 \DRAM_mem_reg[42][22]  ( .D(n7913), .CK(CLK), .QN(n36586) );
  DFF_X1 \DRAM_mem_reg[42][21]  ( .D(n7912), .CK(CLK), .QN(n36584) );
  DFF_X1 \DRAM_mem_reg[42][20]  ( .D(n7911), .CK(CLK), .QN(n36582) );
  DFF_X1 \DRAM_mem_reg[42][19]  ( .D(n7910), .CK(CLK), .QN(n36580) );
  DFF_X1 \DRAM_mem_reg[42][18]  ( .D(n7909), .CK(CLK), .QN(n36578) );
  DFF_X1 \DRAM_mem_reg[42][17]  ( .D(n7908), .CK(CLK), .QN(n36576) );
  DFF_X1 \DRAM_mem_reg[42][16]  ( .D(n7907), .CK(CLK), .QN(n36574) );
  DFF_X1 \DRAM_mem_reg[42][15]  ( .D(n7906), .CK(CLK), .QN(n36572) );
  DFF_X1 \DRAM_mem_reg[42][14]  ( .D(n7905), .CK(CLK), .QN(n36570) );
  DFF_X1 \DRAM_mem_reg[42][13]  ( .D(n7904), .CK(CLK), .QN(n36568) );
  DFF_X1 \DRAM_mem_reg[42][12]  ( .D(n7903), .CK(CLK), .QN(n36566) );
  DFF_X1 \DRAM_mem_reg[42][11]  ( .D(n7902), .CK(CLK), .QN(n36564) );
  DFF_X1 \DRAM_mem_reg[42][10]  ( .D(n7901), .CK(CLK), .QN(n36562) );
  DFF_X1 \DRAM_mem_reg[42][9]  ( .D(n7900), .CK(CLK), .QN(n36560) );
  DFF_X1 \DRAM_mem_reg[42][8]  ( .D(n7899), .CK(CLK), .QN(n36558) );
  DFF_X1 \DRAM_mem_reg[42][7]  ( .D(n7898), .CK(CLK), .QN(n36556) );
  DFF_X1 \DRAM_mem_reg[42][6]  ( .D(n7897), .CK(CLK), .QN(n36554) );
  DFF_X1 \DRAM_mem_reg[42][5]  ( .D(n7896), .CK(CLK), .QN(n36552) );
  DFF_X1 \DRAM_mem_reg[42][4]  ( .D(n7895), .CK(CLK), .QN(n36550) );
  DFF_X1 \DRAM_mem_reg[42][3]  ( .D(n7894), .CK(CLK), .QN(n36548) );
  DFF_X1 \DRAM_mem_reg[42][2]  ( .D(n7893), .CK(CLK), .QN(n36546) );
  DFF_X1 \DRAM_mem_reg[42][1]  ( .D(n7892), .CK(CLK), .QN(n36544) );
  DFF_X1 \DRAM_mem_reg[42][0]  ( .D(n7891), .CK(CLK), .QN(n36542) );
  DFF_X1 \DRAM_mem_reg[43][31]  ( .D(n7890), .CK(CLK), .Q(net253998), .QN(
        n36741) );
  DFF_X1 \DRAM_mem_reg[43][30]  ( .D(n7889), .CK(CLK), .Q(net253997), .QN(
        n36740) );
  DFF_X1 \DRAM_mem_reg[43][29]  ( .D(n7888), .CK(CLK), .Q(net253996), .QN(
        n36739) );
  DFF_X1 \DRAM_mem_reg[43][28]  ( .D(n7887), .CK(CLK), .Q(net253995), .QN(
        n36738) );
  DFF_X1 \DRAM_mem_reg[43][27]  ( .D(n7886), .CK(CLK), .Q(net253994), .QN(
        n36737) );
  DFF_X1 \DRAM_mem_reg[43][26]  ( .D(n7885), .CK(CLK), .Q(net253993), .QN(
        n36736) );
  DFF_X1 \DRAM_mem_reg[43][25]  ( .D(n7884), .CK(CLK), .Q(net253992), .QN(
        n36735) );
  DFF_X1 \DRAM_mem_reg[43][24]  ( .D(n7883), .CK(CLK), .Q(net253991), .QN(
        n36734) );
  DFF_X1 \DRAM_mem_reg[43][23]  ( .D(n7882), .CK(CLK), .Q(net253990), .QN(
        n36949) );
  DFF_X1 \DRAM_mem_reg[43][22]  ( .D(n7881), .CK(CLK), .Q(net253989), .QN(
        n36948) );
  DFF_X1 \DRAM_mem_reg[43][21]  ( .D(n7880), .CK(CLK), .Q(net253988), .QN(
        n36947) );
  DFF_X1 \DRAM_mem_reg[43][20]  ( .D(n7879), .CK(CLK), .Q(net253987), .QN(
        n36946) );
  DFF_X1 \DRAM_mem_reg[43][19]  ( .D(n7878), .CK(CLK), .Q(net253986), .QN(
        n36945) );
  DFF_X1 \DRAM_mem_reg[43][18]  ( .D(n7877), .CK(CLK), .Q(net253985), .QN(
        n36944) );
  DFF_X1 \DRAM_mem_reg[43][17]  ( .D(n7876), .CK(CLK), .Q(net253984), .QN(
        n36943) );
  DFF_X1 \DRAM_mem_reg[43][16]  ( .D(n7875), .CK(CLK), .Q(net253983), .QN(
        n36942) );
  DFF_X1 \DRAM_mem_reg[43][15]  ( .D(n7874), .CK(CLK), .Q(net253982), .QN(
        n36941) );
  DFF_X1 \DRAM_mem_reg[43][14]  ( .D(n7873), .CK(CLK), .Q(net253981), .QN(
        n36940) );
  DFF_X1 \DRAM_mem_reg[43][13]  ( .D(n7872), .CK(CLK), .Q(net253980), .QN(
        n36939) );
  DFF_X1 \DRAM_mem_reg[43][12]  ( .D(n7871), .CK(CLK), .Q(net253979), .QN(
        n36938) );
  DFF_X1 \DRAM_mem_reg[43][11]  ( .D(n7870), .CK(CLK), .Q(net253978), .QN(
        n36937) );
  DFF_X1 \DRAM_mem_reg[43][10]  ( .D(n7869), .CK(CLK), .Q(net253977), .QN(
        n36936) );
  DFF_X1 \DRAM_mem_reg[43][9]  ( .D(n7868), .CK(CLK), .Q(net253976), .QN(
        n36935) );
  DFF_X1 \DRAM_mem_reg[43][8]  ( .D(n7867), .CK(CLK), .Q(net253975), .QN(
        n36934) );
  DFF_X1 \DRAM_mem_reg[43][7]  ( .D(n7866), .CK(CLK), .Q(net253974), .QN(
        n36933) );
  DFF_X1 \DRAM_mem_reg[43][6]  ( .D(n7865), .CK(CLK), .Q(net253973), .QN(
        n36932) );
  DFF_X1 \DRAM_mem_reg[43][5]  ( .D(n7864), .CK(CLK), .Q(net253972), .QN(
        n36931) );
  DFF_X1 \DRAM_mem_reg[43][4]  ( .D(n7863), .CK(CLK), .Q(net253971), .QN(
        n36930) );
  DFF_X1 \DRAM_mem_reg[43][3]  ( .D(n7862), .CK(CLK), .Q(net253970), .QN(
        n36929) );
  DFF_X1 \DRAM_mem_reg[43][2]  ( .D(n7861), .CK(CLK), .Q(net253969), .QN(
        n36928) );
  DFF_X1 \DRAM_mem_reg[43][1]  ( .D(n7860), .CK(CLK), .Q(net253968), .QN(
        n36927) );
  DFF_X1 \DRAM_mem_reg[43][0]  ( .D(n7859), .CK(CLK), .Q(net253967), .QN(
        n36926) );
  DFF_X1 \DRAM_mem_reg[44][31]  ( .D(n7858), .CK(CLK), .QN(n35406) );
  DFF_X1 \DRAM_mem_reg[44][30]  ( .D(n7857), .CK(CLK), .QN(n35397) );
  DFF_X1 \DRAM_mem_reg[44][29]  ( .D(n7856), .CK(CLK), .QN(n35388) );
  DFF_X1 \DRAM_mem_reg[44][28]  ( .D(n7855), .CK(CLK), .QN(n35379) );
  DFF_X1 \DRAM_mem_reg[44][27]  ( .D(n7854), .CK(CLK), .QN(n35370) );
  DFF_X1 \DRAM_mem_reg[44][26]  ( .D(n7853), .CK(CLK), .QN(n35361) );
  DFF_X1 \DRAM_mem_reg[44][25]  ( .D(n7852), .CK(CLK), .QN(n35352) );
  DFF_X1 \DRAM_mem_reg[44][24]  ( .D(n7851), .CK(CLK), .QN(n35343) );
  DFF_X1 \DRAM_mem_reg[44][23]  ( .D(n7850), .CK(CLK), .QN(n35508) );
  DFF_X1 \DRAM_mem_reg[44][22]  ( .D(n7849), .CK(CLK), .QN(n35504) );
  DFF_X1 \DRAM_mem_reg[44][21]  ( .D(n7848), .CK(CLK), .QN(n35500) );
  DFF_X1 \DRAM_mem_reg[44][20]  ( .D(n7847), .CK(CLK), .QN(n35496) );
  DFF_X1 \DRAM_mem_reg[44][19]  ( .D(n7846), .CK(CLK), .QN(n35492) );
  DFF_X1 \DRAM_mem_reg[44][18]  ( .D(n7845), .CK(CLK), .QN(n35488) );
  DFF_X1 \DRAM_mem_reg[44][17]  ( .D(n7844), .CK(CLK), .QN(n35484) );
  DFF_X1 \DRAM_mem_reg[44][16]  ( .D(n7843), .CK(CLK), .QN(n35480) );
  DFF_X1 \DRAM_mem_reg[44][15]  ( .D(n7842), .CK(CLK), .QN(n35476) );
  DFF_X1 \DRAM_mem_reg[44][14]  ( .D(n7841), .CK(CLK), .QN(n35472) );
  DFF_X1 \DRAM_mem_reg[44][13]  ( .D(n7840), .CK(CLK), .QN(n35468) );
  DFF_X1 \DRAM_mem_reg[44][12]  ( .D(n7839), .CK(CLK), .QN(n35464) );
  DFF_X1 \DRAM_mem_reg[44][11]  ( .D(n7838), .CK(CLK), .QN(n35460) );
  DFF_X1 \DRAM_mem_reg[44][10]  ( .D(n7837), .CK(CLK), .QN(n35456) );
  DFF_X1 \DRAM_mem_reg[44][9]  ( .D(n7836), .CK(CLK), .QN(n35452) );
  DFF_X1 \DRAM_mem_reg[44][8]  ( .D(n7835), .CK(CLK), .QN(n35448) );
  DFF_X1 \DRAM_mem_reg[44][7]  ( .D(n7834), .CK(CLK), .QN(n35444) );
  DFF_X1 \DRAM_mem_reg[44][6]  ( .D(n7833), .CK(CLK), .QN(n35440) );
  DFF_X1 \DRAM_mem_reg[44][5]  ( .D(n7832), .CK(CLK), .QN(n35436) );
  DFF_X1 \DRAM_mem_reg[44][4]  ( .D(n7831), .CK(CLK), .QN(n35432) );
  DFF_X1 \DRAM_mem_reg[44][3]  ( .D(n7830), .CK(CLK), .QN(n35428) );
  DFF_X1 \DRAM_mem_reg[44][2]  ( .D(n7829), .CK(CLK), .QN(n35424) );
  DFF_X1 \DRAM_mem_reg[44][1]  ( .D(n7828), .CK(CLK), .QN(n35420) );
  DFF_X1 \DRAM_mem_reg[44][0]  ( .D(n7827), .CK(CLK), .QN(n35416) );
  DFF_X1 \DRAM_mem_reg[45][31]  ( .D(n7826), .CK(CLK), .QN(n35921) );
  DFF_X1 \DRAM_mem_reg[45][30]  ( .D(n7825), .CK(CLK), .QN(n35912) );
  DFF_X1 \DRAM_mem_reg[45][29]  ( .D(n7824), .CK(CLK), .QN(n35903) );
  DFF_X1 \DRAM_mem_reg[45][28]  ( .D(n7823), .CK(CLK), .QN(n35894) );
  DFF_X1 \DRAM_mem_reg[45][27]  ( .D(n7822), .CK(CLK), .QN(n35885) );
  DFF_X1 \DRAM_mem_reg[45][26]  ( .D(n7821), .CK(CLK), .QN(n35876) );
  DFF_X1 \DRAM_mem_reg[45][25]  ( .D(n7820), .CK(CLK), .QN(n35867) );
  DFF_X1 \DRAM_mem_reg[45][24]  ( .D(n7819), .CK(CLK), .QN(n35858) );
  DFF_X1 \DRAM_mem_reg[45][23]  ( .D(n7818), .CK(CLK), .QN(n36172) );
  DFF_X1 \DRAM_mem_reg[45][22]  ( .D(n7817), .CK(CLK), .QN(n36170) );
  DFF_X1 \DRAM_mem_reg[45][21]  ( .D(n7816), .CK(CLK), .QN(n36168) );
  DFF_X1 \DRAM_mem_reg[45][20]  ( .D(n7815), .CK(CLK), .QN(n36166) );
  DFF_X1 \DRAM_mem_reg[45][19]  ( .D(n7814), .CK(CLK), .QN(n36164) );
  DFF_X1 \DRAM_mem_reg[45][18]  ( .D(n7813), .CK(CLK), .QN(n36162) );
  DFF_X1 \DRAM_mem_reg[45][17]  ( .D(n7812), .CK(CLK), .QN(n36160) );
  DFF_X1 \DRAM_mem_reg[45][16]  ( .D(n7811), .CK(CLK), .QN(n36158) );
  DFF_X1 \DRAM_mem_reg[45][15]  ( .D(n7810), .CK(CLK), .QN(n36156) );
  DFF_X1 \DRAM_mem_reg[45][14]  ( .D(n7809), .CK(CLK), .QN(n36154) );
  DFF_X1 \DRAM_mem_reg[45][13]  ( .D(n7808), .CK(CLK), .QN(n36152) );
  DFF_X1 \DRAM_mem_reg[45][12]  ( .D(n7807), .CK(CLK), .QN(n36150) );
  DFF_X1 \DRAM_mem_reg[45][11]  ( .D(n7806), .CK(CLK), .QN(n36148) );
  DFF_X1 \DRAM_mem_reg[45][10]  ( .D(n7805), .CK(CLK), .QN(n36146) );
  DFF_X1 \DRAM_mem_reg[45][9]  ( .D(n7804), .CK(CLK), .QN(n36144) );
  DFF_X1 \DRAM_mem_reg[45][8]  ( .D(n7803), .CK(CLK), .QN(n36142) );
  DFF_X1 \DRAM_mem_reg[45][7]  ( .D(n7802), .CK(CLK), .QN(n36140) );
  DFF_X1 \DRAM_mem_reg[45][6]  ( .D(n7801), .CK(CLK), .QN(n36138) );
  DFF_X1 \DRAM_mem_reg[45][5]  ( .D(n7800), .CK(CLK), .QN(n36136) );
  DFF_X1 \DRAM_mem_reg[45][4]  ( .D(n7799), .CK(CLK), .QN(n36134) );
  DFF_X1 \DRAM_mem_reg[45][3]  ( .D(n7798), .CK(CLK), .QN(n36132) );
  DFF_X1 \DRAM_mem_reg[45][2]  ( .D(n7797), .CK(CLK), .QN(n36130) );
  DFF_X1 \DRAM_mem_reg[45][1]  ( .D(n7796), .CK(CLK), .QN(n36128) );
  DFF_X1 \DRAM_mem_reg[45][0]  ( .D(n7795), .CK(CLK), .QN(n36126) );
  DFF_X1 \DRAM_mem_reg[46][31]  ( .D(n7794), .CK(CLK), .Q(net253966), .QN(
        n37125) );
  DFF_X1 \DRAM_mem_reg[46][30]  ( .D(n7793), .CK(CLK), .Q(net253965), .QN(
        n37124) );
  DFF_X1 \DRAM_mem_reg[46][29]  ( .D(n7792), .CK(CLK), .Q(net253964), .QN(
        n37123) );
  DFF_X1 \DRAM_mem_reg[46][28]  ( .D(n7791), .CK(CLK), .Q(net253963), .QN(
        n37122) );
  DFF_X1 \DRAM_mem_reg[46][27]  ( .D(n7790), .CK(CLK), .Q(net253962), .QN(
        n37121) );
  DFF_X1 \DRAM_mem_reg[46][26]  ( .D(n7789), .CK(CLK), .Q(net253961), .QN(
        n37120) );
  DFF_X1 \DRAM_mem_reg[46][25]  ( .D(n7788), .CK(CLK), .Q(net253960), .QN(
        n37119) );
  DFF_X1 \DRAM_mem_reg[46][24]  ( .D(n7787), .CK(CLK), .Q(net253959), .QN(
        n37118) );
  DFF_X1 \DRAM_mem_reg[46][23]  ( .D(n7786), .CK(CLK), .Q(net253958), .QN(
        n37333) );
  DFF_X1 \DRAM_mem_reg[46][22]  ( .D(n7785), .CK(CLK), .Q(net253957), .QN(
        n37332) );
  DFF_X1 \DRAM_mem_reg[46][21]  ( .D(n7784), .CK(CLK), .Q(net253956), .QN(
        n37331) );
  DFF_X1 \DRAM_mem_reg[46][20]  ( .D(n7783), .CK(CLK), .Q(net253955), .QN(
        n37330) );
  DFF_X1 \DRAM_mem_reg[46][19]  ( .D(n7782), .CK(CLK), .Q(net253954), .QN(
        n37329) );
  DFF_X1 \DRAM_mem_reg[46][18]  ( .D(n7781), .CK(CLK), .Q(net253953), .QN(
        n37328) );
  DFF_X1 \DRAM_mem_reg[46][17]  ( .D(n7780), .CK(CLK), .Q(net253952), .QN(
        n37327) );
  DFF_X1 \DRAM_mem_reg[46][16]  ( .D(n7779), .CK(CLK), .Q(net253951), .QN(
        n37326) );
  DFF_X1 \DRAM_mem_reg[46][15]  ( .D(n7778), .CK(CLK), .Q(net253950), .QN(
        n37325) );
  DFF_X1 \DRAM_mem_reg[46][14]  ( .D(n7777), .CK(CLK), .Q(net253949), .QN(
        n37324) );
  DFF_X1 \DRAM_mem_reg[46][13]  ( .D(n7776), .CK(CLK), .Q(net253948), .QN(
        n37323) );
  DFF_X1 \DRAM_mem_reg[46][12]  ( .D(n7775), .CK(CLK), .Q(net253947), .QN(
        n37322) );
  DFF_X1 \DRAM_mem_reg[46][11]  ( .D(n7774), .CK(CLK), .Q(net253946), .QN(
        n37321) );
  DFF_X1 \DRAM_mem_reg[46][10]  ( .D(n7773), .CK(CLK), .Q(net253945), .QN(
        n37320) );
  DFF_X1 \DRAM_mem_reg[46][9]  ( .D(n7772), .CK(CLK), .Q(net253944), .QN(
        n37319) );
  DFF_X1 \DRAM_mem_reg[46][8]  ( .D(n7771), .CK(CLK), .Q(net253943), .QN(
        n37318) );
  DFF_X1 \DRAM_mem_reg[46][7]  ( .D(n7770), .CK(CLK), .Q(net253942), .QN(
        n37317) );
  DFF_X1 \DRAM_mem_reg[46][6]  ( .D(n7769), .CK(CLK), .Q(net253941), .QN(
        n37316) );
  DFF_X1 \DRAM_mem_reg[46][5]  ( .D(n7768), .CK(CLK), .Q(net253940), .QN(
        n37315) );
  DFF_X1 \DRAM_mem_reg[46][4]  ( .D(n7767), .CK(CLK), .Q(net253939), .QN(
        n37314) );
  DFF_X1 \DRAM_mem_reg[46][3]  ( .D(n7766), .CK(CLK), .Q(net253938), .QN(
        n37313) );
  DFF_X1 \DRAM_mem_reg[46][2]  ( .D(n7765), .CK(CLK), .Q(net253937), .QN(
        n37312) );
  DFF_X1 \DRAM_mem_reg[46][1]  ( .D(n7764), .CK(CLK), .Q(net253936), .QN(
        n37311) );
  DFF_X1 \DRAM_mem_reg[46][0]  ( .D(n7763), .CK(CLK), .Q(net253935), .QN(
        n37310) );
  DFF_X1 \DRAM_mem_reg[47][31]  ( .D(n7762), .CK(CLK), .QN(n36432) );
  DFF_X1 \DRAM_mem_reg[47][30]  ( .D(n7761), .CK(CLK), .QN(n36423) );
  DFF_X1 \DRAM_mem_reg[47][29]  ( .D(n7760), .CK(CLK), .QN(n36414) );
  DFF_X1 \DRAM_mem_reg[47][28]  ( .D(n7759), .CK(CLK), .QN(n36405) );
  DFF_X1 \DRAM_mem_reg[47][27]  ( .D(n7758), .CK(CLK), .QN(n36396) );
  DFF_X1 \DRAM_mem_reg[47][26]  ( .D(n7757), .CK(CLK), .QN(n36387) );
  DFF_X1 \DRAM_mem_reg[47][25]  ( .D(n7756), .CK(CLK), .QN(n36378) );
  DFF_X1 \DRAM_mem_reg[47][24]  ( .D(n7755), .CK(CLK), .QN(n36369) );
  DFF_X1 \DRAM_mem_reg[47][23]  ( .D(n7754), .CK(CLK), .QN(n36636) );
  DFF_X1 \DRAM_mem_reg[47][22]  ( .D(n7753), .CK(CLK), .QN(n36634) );
  DFF_X1 \DRAM_mem_reg[47][21]  ( .D(n7752), .CK(CLK), .QN(n36632) );
  DFF_X1 \DRAM_mem_reg[47][20]  ( .D(n7751), .CK(CLK), .QN(n36630) );
  DFF_X1 \DRAM_mem_reg[47][19]  ( .D(n7750), .CK(CLK), .QN(n36628) );
  DFF_X1 \DRAM_mem_reg[47][18]  ( .D(n7749), .CK(CLK), .QN(n36626) );
  DFF_X1 \DRAM_mem_reg[47][17]  ( .D(n7748), .CK(CLK), .QN(n36624) );
  DFF_X1 \DRAM_mem_reg[47][16]  ( .D(n7747), .CK(CLK), .QN(n36622) );
  DFF_X1 \DRAM_mem_reg[47][15]  ( .D(n7746), .CK(CLK), .QN(n36620) );
  DFF_X1 \DRAM_mem_reg[47][14]  ( .D(n7745), .CK(CLK), .QN(n36618) );
  DFF_X1 \DRAM_mem_reg[47][13]  ( .D(n7744), .CK(CLK), .QN(n36616) );
  DFF_X1 \DRAM_mem_reg[47][12]  ( .D(n7743), .CK(CLK), .QN(n36614) );
  DFF_X1 \DRAM_mem_reg[47][11]  ( .D(n7742), .CK(CLK), .QN(n36612) );
  DFF_X1 \DRAM_mem_reg[47][10]  ( .D(n7741), .CK(CLK), .QN(n36610) );
  DFF_X1 \DRAM_mem_reg[47][9]  ( .D(n7740), .CK(CLK), .QN(n36608) );
  DFF_X1 \DRAM_mem_reg[47][8]  ( .D(n7739), .CK(CLK), .QN(n36606) );
  DFF_X1 \DRAM_mem_reg[47][7]  ( .D(n7738), .CK(CLK), .QN(n36604) );
  DFF_X1 \DRAM_mem_reg[47][6]  ( .D(n7737), .CK(CLK), .QN(n36602) );
  DFF_X1 \DRAM_mem_reg[47][5]  ( .D(n7736), .CK(CLK), .QN(n36600) );
  DFF_X1 \DRAM_mem_reg[47][4]  ( .D(n7735), .CK(CLK), .QN(n36598) );
  DFF_X1 \DRAM_mem_reg[47][3]  ( .D(n7734), .CK(CLK), .QN(n36596) );
  DFF_X1 \DRAM_mem_reg[47][2]  ( .D(n7733), .CK(CLK), .QN(n36594) );
  DFF_X1 \DRAM_mem_reg[47][1]  ( .D(n7732), .CK(CLK), .QN(n36592) );
  DFF_X1 \DRAM_mem_reg[47][0]  ( .D(n7731), .CK(CLK), .QN(n36590) );
  DFF_X1 \DRAM_mem_reg[48][31]  ( .D(n7730), .CK(CLK), .QN(n35685) );
  DFF_X1 \DRAM_mem_reg[48][30]  ( .D(n7729), .CK(CLK), .QN(n35684) );
  DFF_X1 \DRAM_mem_reg[48][29]  ( .D(n7728), .CK(CLK), .QN(n35683) );
  DFF_X1 \DRAM_mem_reg[48][28]  ( .D(n7727), .CK(CLK), .QN(n35682) );
  DFF_X1 \DRAM_mem_reg[48][27]  ( .D(n7726), .CK(CLK), .QN(n35681) );
  DFF_X1 \DRAM_mem_reg[48][26]  ( .D(n7725), .CK(CLK), .QN(n35680) );
  DFF_X1 \DRAM_mem_reg[48][25]  ( .D(n7724), .CK(CLK), .QN(n35679) );
  DFF_X1 \DRAM_mem_reg[48][24]  ( .D(n7723), .CK(CLK), .QN(n35678) );
  DFF_X1 \DRAM_mem_reg[48][23]  ( .D(n7722), .CK(CLK), .QN(n35781) );
  DFF_X1 \DRAM_mem_reg[48][22]  ( .D(n7721), .CK(CLK), .QN(n35780) );
  DFF_X1 \DRAM_mem_reg[48][21]  ( .D(n7720), .CK(CLK), .QN(n35779) );
  DFF_X1 \DRAM_mem_reg[48][20]  ( .D(n7719), .CK(CLK), .QN(n35778) );
  DFF_X1 \DRAM_mem_reg[48][19]  ( .D(n7718), .CK(CLK), .QN(n35777) );
  DFF_X1 \DRAM_mem_reg[48][18]  ( .D(n7717), .CK(CLK), .QN(n35776) );
  DFF_X1 \DRAM_mem_reg[48][17]  ( .D(n7716), .CK(CLK), .QN(n35775) );
  DFF_X1 \DRAM_mem_reg[48][16]  ( .D(n7715), .CK(CLK), .QN(n35774) );
  DFF_X1 \DRAM_mem_reg[48][15]  ( .D(n7714), .CK(CLK), .QN(n35773) );
  DFF_X1 \DRAM_mem_reg[48][14]  ( .D(n7713), .CK(CLK), .QN(n35772) );
  DFF_X1 \DRAM_mem_reg[48][13]  ( .D(n7712), .CK(CLK), .QN(n35771) );
  DFF_X1 \DRAM_mem_reg[48][12]  ( .D(n7711), .CK(CLK), .QN(n35770) );
  DFF_X1 \DRAM_mem_reg[48][11]  ( .D(n7710), .CK(CLK), .QN(n35769) );
  DFF_X1 \DRAM_mem_reg[48][10]  ( .D(n7709), .CK(CLK), .QN(n35768) );
  DFF_X1 \DRAM_mem_reg[48][9]  ( .D(n7708), .CK(CLK), .QN(n35767) );
  DFF_X1 \DRAM_mem_reg[48][8]  ( .D(n7707), .CK(CLK), .QN(n35766) );
  DFF_X1 \DRAM_mem_reg[48][7]  ( .D(n7706), .CK(CLK), .QN(n35765) );
  DFF_X1 \DRAM_mem_reg[48][6]  ( .D(n7705), .CK(CLK), .QN(n35764) );
  DFF_X1 \DRAM_mem_reg[48][5]  ( .D(n7704), .CK(CLK), .QN(n35763) );
  DFF_X1 \DRAM_mem_reg[48][4]  ( .D(n7703), .CK(CLK), .QN(n35762) );
  DFF_X1 \DRAM_mem_reg[48][3]  ( .D(n7702), .CK(CLK), .QN(n35761) );
  DFF_X1 \DRAM_mem_reg[48][2]  ( .D(n7701), .CK(CLK), .QN(n35760) );
  DFF_X1 \DRAM_mem_reg[48][1]  ( .D(n7700), .CK(CLK), .QN(n35759) );
  DFF_X1 \DRAM_mem_reg[48][0]  ( .D(n7699), .CK(CLK), .QN(n35758) );
  DFF_X1 \DRAM_mem_reg[49][31]  ( .D(n7698), .CK(CLK), .Q(net253934), .QN(
        n37117) );
  DFF_X1 \DRAM_mem_reg[49][30]  ( .D(n7697), .CK(CLK), .Q(net253933), .QN(
        n37116) );
  DFF_X1 \DRAM_mem_reg[49][29]  ( .D(n7696), .CK(CLK), .Q(net253932), .QN(
        n37115) );
  DFF_X1 \DRAM_mem_reg[49][28]  ( .D(n7695), .CK(CLK), .Q(net253931), .QN(
        n37114) );
  DFF_X1 \DRAM_mem_reg[49][27]  ( .D(n7694), .CK(CLK), .Q(net253930), .QN(
        n37113) );
  DFF_X1 \DRAM_mem_reg[49][26]  ( .D(n7693), .CK(CLK), .Q(net253929), .QN(
        n37112) );
  DFF_X1 \DRAM_mem_reg[49][25]  ( .D(n7692), .CK(CLK), .Q(net253928), .QN(
        n37111) );
  DFF_X1 \DRAM_mem_reg[49][24]  ( .D(n7691), .CK(CLK), .Q(net253927), .QN(
        n37110) );
  DFF_X1 \DRAM_mem_reg[49][23]  ( .D(n7690), .CK(CLK), .Q(net253926), .QN(
        n37309) );
  DFF_X1 \DRAM_mem_reg[49][22]  ( .D(n7689), .CK(CLK), .Q(net253925), .QN(
        n37308) );
  DFF_X1 \DRAM_mem_reg[49][21]  ( .D(n7688), .CK(CLK), .Q(net253924), .QN(
        n37307) );
  DFF_X1 \DRAM_mem_reg[49][20]  ( .D(n7687), .CK(CLK), .Q(net253923), .QN(
        n37306) );
  DFF_X1 \DRAM_mem_reg[49][19]  ( .D(n7686), .CK(CLK), .Q(net253922), .QN(
        n37305) );
  DFF_X1 \DRAM_mem_reg[49][18]  ( .D(n7685), .CK(CLK), .Q(net253921), .QN(
        n37304) );
  DFF_X1 \DRAM_mem_reg[49][17]  ( .D(n7684), .CK(CLK), .Q(net253920), .QN(
        n37303) );
  DFF_X1 \DRAM_mem_reg[49][16]  ( .D(n7683), .CK(CLK), .Q(net253919), .QN(
        n37302) );
  DFF_X1 \DRAM_mem_reg[49][15]  ( .D(n7682), .CK(CLK), .Q(net253918), .QN(
        n37301) );
  DFF_X1 \DRAM_mem_reg[49][14]  ( .D(n7681), .CK(CLK), .Q(net253917), .QN(
        n37300) );
  DFF_X1 \DRAM_mem_reg[49][13]  ( .D(n7680), .CK(CLK), .Q(net253916), .QN(
        n37299) );
  DFF_X1 \DRAM_mem_reg[49][12]  ( .D(n7679), .CK(CLK), .Q(net253915), .QN(
        n37298) );
  DFF_X1 \DRAM_mem_reg[49][11]  ( .D(n7678), .CK(CLK), .Q(net253914), .QN(
        n37297) );
  DFF_X1 \DRAM_mem_reg[49][10]  ( .D(n7677), .CK(CLK), .Q(net253913), .QN(
        n37296) );
  DFF_X1 \DRAM_mem_reg[49][9]  ( .D(n7676), .CK(CLK), .Q(net253912), .QN(
        n37295) );
  DFF_X1 \DRAM_mem_reg[49][8]  ( .D(n7675), .CK(CLK), .Q(net253911), .QN(
        n37294) );
  DFF_X1 \DRAM_mem_reg[49][7]  ( .D(n7674), .CK(CLK), .Q(net253910), .QN(
        n37293) );
  DFF_X1 \DRAM_mem_reg[49][6]  ( .D(n7673), .CK(CLK), .Q(net253909), .QN(
        n37292) );
  DFF_X1 \DRAM_mem_reg[49][5]  ( .D(n7672), .CK(CLK), .Q(net253908), .QN(
        n37291) );
  DFF_X1 \DRAM_mem_reg[49][4]  ( .D(n7671), .CK(CLK), .Q(net253907), .QN(
        n37290) );
  DFF_X1 \DRAM_mem_reg[49][3]  ( .D(n7670), .CK(CLK), .Q(net253906), .QN(
        n37289) );
  DFF_X1 \DRAM_mem_reg[49][2]  ( .D(n7669), .CK(CLK), .Q(net253905), .QN(
        n37288) );
  DFF_X1 \DRAM_mem_reg[49][1]  ( .D(n7668), .CK(CLK), .Q(net253904), .QN(
        n37287) );
  DFF_X1 \DRAM_mem_reg[49][0]  ( .D(n7667), .CK(CLK), .Q(net253903), .QN(
        n37286) );
  DFF_X1 \DRAM_mem_reg[50][31]  ( .D(n7666), .CK(CLK), .QN(n36197) );
  DFF_X1 \DRAM_mem_reg[50][30]  ( .D(n7665), .CK(CLK), .QN(n36196) );
  DFF_X1 \DRAM_mem_reg[50][29]  ( .D(n7664), .CK(CLK), .QN(n36195) );
  DFF_X1 \DRAM_mem_reg[50][28]  ( .D(n7663), .CK(CLK), .QN(n36194) );
  DFF_X1 \DRAM_mem_reg[50][27]  ( .D(n7662), .CK(CLK), .QN(n36193) );
  DFF_X1 \DRAM_mem_reg[50][26]  ( .D(n7661), .CK(CLK), .QN(n36192) );
  DFF_X1 \DRAM_mem_reg[50][25]  ( .D(n7660), .CK(CLK), .QN(n36191) );
  DFF_X1 \DRAM_mem_reg[50][24]  ( .D(n7659), .CK(CLK), .QN(n36190) );
  DFF_X1 \DRAM_mem_reg[50][23]  ( .D(n7658), .CK(CLK), .QN(n36293) );
  DFF_X1 \DRAM_mem_reg[50][22]  ( .D(n7657), .CK(CLK), .QN(n36292) );
  DFF_X1 \DRAM_mem_reg[50][21]  ( .D(n7656), .CK(CLK), .QN(n36291) );
  DFF_X1 \DRAM_mem_reg[50][20]  ( .D(n7655), .CK(CLK), .QN(n36290) );
  DFF_X1 \DRAM_mem_reg[50][19]  ( .D(n7654), .CK(CLK), .QN(n36289) );
  DFF_X1 \DRAM_mem_reg[50][18]  ( .D(n7653), .CK(CLK), .QN(n36288) );
  DFF_X1 \DRAM_mem_reg[50][17]  ( .D(n7652), .CK(CLK), .QN(n36287) );
  DFF_X1 \DRAM_mem_reg[50][16]  ( .D(n7651), .CK(CLK), .QN(n36286) );
  DFF_X1 \DRAM_mem_reg[50][15]  ( .D(n7650), .CK(CLK), .QN(n36285) );
  DFF_X1 \DRAM_mem_reg[50][14]  ( .D(n7649), .CK(CLK), .QN(n36284) );
  DFF_X1 \DRAM_mem_reg[50][13]  ( .D(n7648), .CK(CLK), .QN(n36283) );
  DFF_X1 \DRAM_mem_reg[50][12]  ( .D(n7647), .CK(CLK), .QN(n36282) );
  DFF_X1 \DRAM_mem_reg[50][11]  ( .D(n7646), .CK(CLK), .QN(n36281) );
  DFF_X1 \DRAM_mem_reg[50][10]  ( .D(n7645), .CK(CLK), .QN(n36280) );
  DFF_X1 \DRAM_mem_reg[50][9]  ( .D(n7644), .CK(CLK), .QN(n36279) );
  DFF_X1 \DRAM_mem_reg[50][8]  ( .D(n7643), .CK(CLK), .QN(n36278) );
  DFF_X1 \DRAM_mem_reg[50][7]  ( .D(n7642), .CK(CLK), .QN(n36277) );
  DFF_X1 \DRAM_mem_reg[50][6]  ( .D(n7641), .CK(CLK), .QN(n36276) );
  DFF_X1 \DRAM_mem_reg[50][5]  ( .D(n7640), .CK(CLK), .QN(n36275) );
  DFF_X1 \DRAM_mem_reg[50][4]  ( .D(n7639), .CK(CLK), .QN(n36274) );
  DFF_X1 \DRAM_mem_reg[50][3]  ( .D(n7638), .CK(CLK), .QN(n36273) );
  DFF_X1 \DRAM_mem_reg[50][2]  ( .D(n7637), .CK(CLK), .QN(n36272) );
  DFF_X1 \DRAM_mem_reg[50][1]  ( .D(n7636), .CK(CLK), .QN(n36271) );
  DFF_X1 \DRAM_mem_reg[50][0]  ( .D(n7635), .CK(CLK), .QN(n36270) );
  DFF_X1 \DRAM_mem_reg[51][31]  ( .D(n7634), .CK(CLK), .Q(net253902), .QN(
        n36733) );
  DFF_X1 \DRAM_mem_reg[51][30]  ( .D(n7633), .CK(CLK), .Q(net253901), .QN(
        n36732) );
  DFF_X1 \DRAM_mem_reg[51][29]  ( .D(n7632), .CK(CLK), .Q(net253900), .QN(
        n36731) );
  DFF_X1 \DRAM_mem_reg[51][28]  ( .D(n7631), .CK(CLK), .Q(net253899), .QN(
        n36730) );
  DFF_X1 \DRAM_mem_reg[51][27]  ( .D(n7630), .CK(CLK), .Q(net253898), .QN(
        n36729) );
  DFF_X1 \DRAM_mem_reg[51][26]  ( .D(n7629), .CK(CLK), .Q(net253897), .QN(
        n36728) );
  DFF_X1 \DRAM_mem_reg[51][25]  ( .D(n7628), .CK(CLK), .Q(net253896), .QN(
        n36727) );
  DFF_X1 \DRAM_mem_reg[51][24]  ( .D(n7627), .CK(CLK), .Q(net253895), .QN(
        n36726) );
  DFF_X1 \DRAM_mem_reg[51][23]  ( .D(n7626), .CK(CLK), .Q(net253894), .QN(
        n36925) );
  DFF_X1 \DRAM_mem_reg[51][22]  ( .D(n7625), .CK(CLK), .Q(net253893), .QN(
        n36924) );
  DFF_X1 \DRAM_mem_reg[51][21]  ( .D(n7624), .CK(CLK), .Q(net253892), .QN(
        n36923) );
  DFF_X1 \DRAM_mem_reg[51][20]  ( .D(n7623), .CK(CLK), .Q(net253891), .QN(
        n36922) );
  DFF_X1 \DRAM_mem_reg[51][19]  ( .D(n7622), .CK(CLK), .Q(net253890), .QN(
        n36921) );
  DFF_X1 \DRAM_mem_reg[51][18]  ( .D(n7621), .CK(CLK), .Q(net253889), .QN(
        n36920) );
  DFF_X1 \DRAM_mem_reg[51][17]  ( .D(n7620), .CK(CLK), .Q(net253888), .QN(
        n36919) );
  DFF_X1 \DRAM_mem_reg[51][16]  ( .D(n7619), .CK(CLK), .Q(net253887), .QN(
        n36918) );
  DFF_X1 \DRAM_mem_reg[51][15]  ( .D(n7618), .CK(CLK), .Q(net253886), .QN(
        n36917) );
  DFF_X1 \DRAM_mem_reg[51][14]  ( .D(n7617), .CK(CLK), .Q(net253885), .QN(
        n36916) );
  DFF_X1 \DRAM_mem_reg[51][13]  ( .D(n7616), .CK(CLK), .Q(net253884), .QN(
        n36915) );
  DFF_X1 \DRAM_mem_reg[51][12]  ( .D(n7615), .CK(CLK), .Q(net253883), .QN(
        n36914) );
  DFF_X1 \DRAM_mem_reg[51][11]  ( .D(n7614), .CK(CLK), .Q(net253882), .QN(
        n36913) );
  DFF_X1 \DRAM_mem_reg[51][10]  ( .D(n7613), .CK(CLK), .Q(net253881), .QN(
        n36912) );
  DFF_X1 \DRAM_mem_reg[51][9]  ( .D(n7612), .CK(CLK), .Q(net253880), .QN(
        n36911) );
  DFF_X1 \DRAM_mem_reg[51][8]  ( .D(n7611), .CK(CLK), .Q(net253879), .QN(
        n36910) );
  DFF_X1 \DRAM_mem_reg[51][7]  ( .D(n7610), .CK(CLK), .Q(net253878), .QN(
        n36909) );
  DFF_X1 \DRAM_mem_reg[51][6]  ( .D(n7609), .CK(CLK), .Q(net253877), .QN(
        n36908) );
  DFF_X1 \DRAM_mem_reg[51][5]  ( .D(n7608), .CK(CLK), .Q(net253876), .QN(
        n36907) );
  DFF_X1 \DRAM_mem_reg[51][4]  ( .D(n7607), .CK(CLK), .Q(net253875), .QN(
        n36906) );
  DFF_X1 \DRAM_mem_reg[51][3]  ( .D(n7606), .CK(CLK), .Q(net253874), .QN(
        n36905) );
  DFF_X1 \DRAM_mem_reg[51][2]  ( .D(n7605), .CK(CLK), .Q(net253873), .QN(
        n36904) );
  DFF_X1 \DRAM_mem_reg[51][1]  ( .D(n7604), .CK(CLK), .Q(net253872), .QN(
        n36903) );
  DFF_X1 \DRAM_mem_reg[51][0]  ( .D(n7603), .CK(CLK), .Q(net253871), .QN(
        n36902) );
  DFF_X1 \DRAM_mem_reg[52][31]  ( .D(n7602), .CK(CLK), .QN(n35411) );
  DFF_X1 \DRAM_mem_reg[52][30]  ( .D(n7601), .CK(CLK), .QN(n35402) );
  DFF_X1 \DRAM_mem_reg[52][29]  ( .D(n7600), .CK(CLK), .QN(n35393) );
  DFF_X1 \DRAM_mem_reg[52][28]  ( .D(n7599), .CK(CLK), .QN(n35384) );
  DFF_X1 \DRAM_mem_reg[52][27]  ( .D(n7598), .CK(CLK), .QN(n35375) );
  DFF_X1 \DRAM_mem_reg[52][26]  ( .D(n7597), .CK(CLK), .QN(n35366) );
  DFF_X1 \DRAM_mem_reg[52][25]  ( .D(n7596), .CK(CLK), .QN(n35357) );
  DFF_X1 \DRAM_mem_reg[52][24]  ( .D(n7595), .CK(CLK), .QN(n35348) );
  DFF_X1 \DRAM_mem_reg[52][23]  ( .D(n7594), .CK(CLK), .QN(n35565) );
  DFF_X1 \DRAM_mem_reg[52][22]  ( .D(n7593), .CK(CLK), .QN(n35563) );
  DFF_X1 \DRAM_mem_reg[52][21]  ( .D(n7592), .CK(CLK), .QN(n35561) );
  DFF_X1 \DRAM_mem_reg[52][20]  ( .D(n7591), .CK(CLK), .QN(n35559) );
  DFF_X1 \DRAM_mem_reg[52][19]  ( .D(n7590), .CK(CLK), .QN(n35557) );
  DFF_X1 \DRAM_mem_reg[52][18]  ( .D(n7589), .CK(CLK), .QN(n35555) );
  DFF_X1 \DRAM_mem_reg[52][17]  ( .D(n7588), .CK(CLK), .QN(n35553) );
  DFF_X1 \DRAM_mem_reg[52][16]  ( .D(n7587), .CK(CLK), .QN(n35551) );
  DFF_X1 \DRAM_mem_reg[52][15]  ( .D(n7586), .CK(CLK), .QN(n35549) );
  DFF_X1 \DRAM_mem_reg[52][14]  ( .D(n7585), .CK(CLK), .QN(n35547) );
  DFF_X1 \DRAM_mem_reg[52][13]  ( .D(n7584), .CK(CLK), .QN(n35545) );
  DFF_X1 \DRAM_mem_reg[52][12]  ( .D(n7583), .CK(CLK), .QN(n35543) );
  DFF_X1 \DRAM_mem_reg[52][11]  ( .D(n7582), .CK(CLK), .QN(n35541) );
  DFF_X1 \DRAM_mem_reg[52][10]  ( .D(n7581), .CK(CLK), .QN(n35539) );
  DFF_X1 \DRAM_mem_reg[52][9]  ( .D(n7580), .CK(CLK), .QN(n35537) );
  DFF_X1 \DRAM_mem_reg[52][8]  ( .D(n7579), .CK(CLK), .QN(n35535) );
  DFF_X1 \DRAM_mem_reg[52][7]  ( .D(n7578), .CK(CLK), .QN(n35533) );
  DFF_X1 \DRAM_mem_reg[52][6]  ( .D(n7577), .CK(CLK), .QN(n35531) );
  DFF_X1 \DRAM_mem_reg[52][5]  ( .D(n7576), .CK(CLK), .QN(n35529) );
  DFF_X1 \DRAM_mem_reg[52][4]  ( .D(n7575), .CK(CLK), .QN(n35527) );
  DFF_X1 \DRAM_mem_reg[52][3]  ( .D(n7574), .CK(CLK), .QN(n35525) );
  DFF_X1 \DRAM_mem_reg[52][2]  ( .D(n7573), .CK(CLK), .QN(n35523) );
  DFF_X1 \DRAM_mem_reg[52][1]  ( .D(n7572), .CK(CLK), .QN(n35521) );
  DFF_X1 \DRAM_mem_reg[52][0]  ( .D(n7571), .CK(CLK), .QN(n35519) );
  DFF_X1 \DRAM_mem_reg[53][31]  ( .D(n7570), .CK(CLK), .QN(n35922) );
  DFF_X1 \DRAM_mem_reg[53][30]  ( .D(n7569), .CK(CLK), .QN(n35913) );
  DFF_X1 \DRAM_mem_reg[53][29]  ( .D(n7568), .CK(CLK), .QN(n35904) );
  DFF_X1 \DRAM_mem_reg[53][28]  ( .D(n7567), .CK(CLK), .QN(n35895) );
  DFF_X1 \DRAM_mem_reg[53][27]  ( .D(n7566), .CK(CLK), .QN(n35886) );
  DFF_X1 \DRAM_mem_reg[53][26]  ( .D(n7565), .CK(CLK), .QN(n35877) );
  DFF_X1 \DRAM_mem_reg[53][25]  ( .D(n7564), .CK(CLK), .QN(n35868) );
  DFF_X1 \DRAM_mem_reg[53][24]  ( .D(n7563), .CK(CLK), .QN(n35859) );
  DFF_X1 \DRAM_mem_reg[53][23]  ( .D(n7562), .CK(CLK), .QN(n36021) );
  DFF_X1 \DRAM_mem_reg[53][22]  ( .D(n7561), .CK(CLK), .QN(n36017) );
  DFF_X1 \DRAM_mem_reg[53][21]  ( .D(n7560), .CK(CLK), .QN(n36013) );
  DFF_X1 \DRAM_mem_reg[53][20]  ( .D(n7559), .CK(CLK), .QN(n36009) );
  DFF_X1 \DRAM_mem_reg[53][19]  ( .D(n7558), .CK(CLK), .QN(n36005) );
  DFF_X1 \DRAM_mem_reg[53][18]  ( .D(n7557), .CK(CLK), .QN(n36001) );
  DFF_X1 \DRAM_mem_reg[53][17]  ( .D(n7556), .CK(CLK), .QN(n35997) );
  DFF_X1 \DRAM_mem_reg[53][16]  ( .D(n7555), .CK(CLK), .QN(n35993) );
  DFF_X1 \DRAM_mem_reg[53][15]  ( .D(n7554), .CK(CLK), .QN(n35989) );
  DFF_X1 \DRAM_mem_reg[53][14]  ( .D(n7553), .CK(CLK), .QN(n35985) );
  DFF_X1 \DRAM_mem_reg[53][13]  ( .D(n7552), .CK(CLK), .QN(n35981) );
  DFF_X1 \DRAM_mem_reg[53][12]  ( .D(n7551), .CK(CLK), .QN(n35977) );
  DFF_X1 \DRAM_mem_reg[53][11]  ( .D(n7550), .CK(CLK), .QN(n35973) );
  DFF_X1 \DRAM_mem_reg[53][10]  ( .D(n7549), .CK(CLK), .QN(n35969) );
  DFF_X1 \DRAM_mem_reg[53][9]  ( .D(n7548), .CK(CLK), .QN(n35965) );
  DFF_X1 \DRAM_mem_reg[53][8]  ( .D(n7547), .CK(CLK), .QN(n35961) );
  DFF_X1 \DRAM_mem_reg[53][7]  ( .D(n7546), .CK(CLK), .QN(n35957) );
  DFF_X1 \DRAM_mem_reg[53][6]  ( .D(n7545), .CK(CLK), .QN(n35953) );
  DFF_X1 \DRAM_mem_reg[53][5]  ( .D(n7544), .CK(CLK), .QN(n35949) );
  DFF_X1 \DRAM_mem_reg[53][4]  ( .D(n7543), .CK(CLK), .QN(n35945) );
  DFF_X1 \DRAM_mem_reg[53][3]  ( .D(n7542), .CK(CLK), .QN(n35941) );
  DFF_X1 \DRAM_mem_reg[53][2]  ( .D(n7541), .CK(CLK), .QN(n35937) );
  DFF_X1 \DRAM_mem_reg[53][1]  ( .D(n7540), .CK(CLK), .QN(n35933) );
  DFF_X1 \DRAM_mem_reg[53][0]  ( .D(n7539), .CK(CLK), .QN(n35929) );
  DFF_X1 \DRAM_mem_reg[54][31]  ( .D(n7538), .CK(CLK), .Q(net253870), .QN(
        n37109) );
  DFF_X1 \DRAM_mem_reg[54][30]  ( .D(n7537), .CK(CLK), .Q(net253869), .QN(
        n37108) );
  DFF_X1 \DRAM_mem_reg[54][29]  ( .D(n7536), .CK(CLK), .Q(net253868), .QN(
        n37107) );
  DFF_X1 \DRAM_mem_reg[54][28]  ( .D(n7535), .CK(CLK), .Q(net253867), .QN(
        n37106) );
  DFF_X1 \DRAM_mem_reg[54][27]  ( .D(n7534), .CK(CLK), .Q(net253866), .QN(
        n37105) );
  DFF_X1 \DRAM_mem_reg[54][26]  ( .D(n7533), .CK(CLK), .Q(net253865), .QN(
        n37104) );
  DFF_X1 \DRAM_mem_reg[54][25]  ( .D(n7532), .CK(CLK), .Q(net253864), .QN(
        n37103) );
  DFF_X1 \DRAM_mem_reg[54][24]  ( .D(n7531), .CK(CLK), .Q(net253863), .QN(
        n37102) );
  DFF_X1 \DRAM_mem_reg[54][23]  ( .D(n7530), .CK(CLK), .Q(net253862), .QN(
        n37285) );
  DFF_X1 \DRAM_mem_reg[54][22]  ( .D(n7529), .CK(CLK), .Q(net253861), .QN(
        n37284) );
  DFF_X1 \DRAM_mem_reg[54][21]  ( .D(n7528), .CK(CLK), .Q(net253860), .QN(
        n37283) );
  DFF_X1 \DRAM_mem_reg[54][20]  ( .D(n7527), .CK(CLK), .Q(net253859), .QN(
        n37282) );
  DFF_X1 \DRAM_mem_reg[54][19]  ( .D(n7526), .CK(CLK), .Q(net253858), .QN(
        n37281) );
  DFF_X1 \DRAM_mem_reg[54][18]  ( .D(n7525), .CK(CLK), .Q(net253857), .QN(
        n37280) );
  DFF_X1 \DRAM_mem_reg[54][17]  ( .D(n7524), .CK(CLK), .Q(net253856), .QN(
        n37279) );
  DFF_X1 \DRAM_mem_reg[54][16]  ( .D(n7523), .CK(CLK), .Q(net253855), .QN(
        n37278) );
  DFF_X1 \DRAM_mem_reg[54][15]  ( .D(n7522), .CK(CLK), .Q(net253854), .QN(
        n37277) );
  DFF_X1 \DRAM_mem_reg[54][14]  ( .D(n7521), .CK(CLK), .Q(net253853), .QN(
        n37276) );
  DFF_X1 \DRAM_mem_reg[54][13]  ( .D(n7520), .CK(CLK), .Q(net253852), .QN(
        n37275) );
  DFF_X1 \DRAM_mem_reg[54][12]  ( .D(n7519), .CK(CLK), .Q(net253851), .QN(
        n37274) );
  DFF_X1 \DRAM_mem_reg[54][11]  ( .D(n7518), .CK(CLK), .Q(net253850), .QN(
        n37273) );
  DFF_X1 \DRAM_mem_reg[54][10]  ( .D(n7517), .CK(CLK), .Q(net253849), .QN(
        n37272) );
  DFF_X1 \DRAM_mem_reg[54][9]  ( .D(n7516), .CK(CLK), .Q(net253848), .QN(
        n37271) );
  DFF_X1 \DRAM_mem_reg[54][8]  ( .D(n7515), .CK(CLK), .Q(net253847), .QN(
        n37270) );
  DFF_X1 \DRAM_mem_reg[54][7]  ( .D(n7514), .CK(CLK), .Q(net253846), .QN(
        n37269) );
  DFF_X1 \DRAM_mem_reg[54][6]  ( .D(n7513), .CK(CLK), .Q(net253845), .QN(
        n37268) );
  DFF_X1 \DRAM_mem_reg[54][5]  ( .D(n7512), .CK(CLK), .Q(net253844), .QN(
        n37267) );
  DFF_X1 \DRAM_mem_reg[54][4]  ( .D(n7511), .CK(CLK), .Q(net253843), .QN(
        n37266) );
  DFF_X1 \DRAM_mem_reg[54][3]  ( .D(n7510), .CK(CLK), .Q(net253842), .QN(
        n37265) );
  DFF_X1 \DRAM_mem_reg[54][2]  ( .D(n7509), .CK(CLK), .Q(net253841), .QN(
        n37264) );
  DFF_X1 \DRAM_mem_reg[54][1]  ( .D(n7508), .CK(CLK), .Q(net253840), .QN(
        n37263) );
  DFF_X1 \DRAM_mem_reg[54][0]  ( .D(n7507), .CK(CLK), .Q(net253839), .QN(
        n37262) );
  DFF_X1 \DRAM_mem_reg[55][31]  ( .D(n7506), .CK(CLK), .QN(n36437) );
  DFF_X1 \DRAM_mem_reg[55][30]  ( .D(n7505), .CK(CLK), .QN(n36428) );
  DFF_X1 \DRAM_mem_reg[55][29]  ( .D(n7504), .CK(CLK), .QN(n36419) );
  DFF_X1 \DRAM_mem_reg[55][28]  ( .D(n7503), .CK(CLK), .QN(n36410) );
  DFF_X1 \DRAM_mem_reg[55][27]  ( .D(n7502), .CK(CLK), .QN(n36401) );
  DFF_X1 \DRAM_mem_reg[55][26]  ( .D(n7501), .CK(CLK), .QN(n36392) );
  DFF_X1 \DRAM_mem_reg[55][25]  ( .D(n7500), .CK(CLK), .QN(n36383) );
  DFF_X1 \DRAM_mem_reg[55][24]  ( .D(n7499), .CK(CLK), .QN(n36374) );
  DFF_X1 \DRAM_mem_reg[55][23]  ( .D(n7498), .CK(CLK), .QN(n36685) );
  DFF_X1 \DRAM_mem_reg[55][22]  ( .D(n7497), .CK(CLK), .QN(n36683) );
  DFF_X1 \DRAM_mem_reg[55][21]  ( .D(n7496), .CK(CLK), .QN(n36681) );
  DFF_X1 \DRAM_mem_reg[55][20]  ( .D(n7495), .CK(CLK), .QN(n36679) );
  DFF_X1 \DRAM_mem_reg[55][19]  ( .D(n7494), .CK(CLK), .QN(n36677) );
  DFF_X1 \DRAM_mem_reg[55][18]  ( .D(n7493), .CK(CLK), .QN(n36675) );
  DFF_X1 \DRAM_mem_reg[55][17]  ( .D(n7492), .CK(CLK), .QN(n36673) );
  DFF_X1 \DRAM_mem_reg[55][16]  ( .D(n7491), .CK(CLK), .QN(n36671) );
  DFF_X1 \DRAM_mem_reg[55][15]  ( .D(n7490), .CK(CLK), .QN(n36669) );
  DFF_X1 \DRAM_mem_reg[55][14]  ( .D(n7489), .CK(CLK), .QN(n36667) );
  DFF_X1 \DRAM_mem_reg[55][13]  ( .D(n7488), .CK(CLK), .QN(n36665) );
  DFF_X1 \DRAM_mem_reg[55][12]  ( .D(n7487), .CK(CLK), .QN(n36663) );
  DFF_X1 \DRAM_mem_reg[55][11]  ( .D(n7486), .CK(CLK), .QN(n36661) );
  DFF_X1 \DRAM_mem_reg[55][10]  ( .D(n7485), .CK(CLK), .QN(n36659) );
  DFF_X1 \DRAM_mem_reg[55][9]  ( .D(n7484), .CK(CLK), .QN(n36657) );
  DFF_X1 \DRAM_mem_reg[55][8]  ( .D(n7483), .CK(CLK), .QN(n36655) );
  DFF_X1 \DRAM_mem_reg[55][7]  ( .D(n7482), .CK(CLK), .QN(n36653) );
  DFF_X1 \DRAM_mem_reg[55][6]  ( .D(n7481), .CK(CLK), .QN(n36651) );
  DFF_X1 \DRAM_mem_reg[55][5]  ( .D(n7480), .CK(CLK), .QN(n36649) );
  DFF_X1 \DRAM_mem_reg[55][4]  ( .D(n7479), .CK(CLK), .QN(n36647) );
  DFF_X1 \DRAM_mem_reg[55][3]  ( .D(n7478), .CK(CLK), .QN(n36645) );
  DFF_X1 \DRAM_mem_reg[55][2]  ( .D(n7477), .CK(CLK), .QN(n36643) );
  DFF_X1 \DRAM_mem_reg[55][1]  ( .D(n7476), .CK(CLK), .QN(n36641) );
  DFF_X1 \DRAM_mem_reg[55][0]  ( .D(n7475), .CK(CLK), .QN(n36639) );
  DFF_X1 \DRAM_mem_reg[56][31]  ( .D(n7474), .CK(CLK), .Q(net253838), .QN(
        n36725) );
  DFF_X1 \DRAM_mem_reg[56][30]  ( .D(n7473), .CK(CLK), .Q(net253837), .QN(
        n36724) );
  DFF_X1 \DRAM_mem_reg[56][29]  ( .D(n7472), .CK(CLK), .Q(net253836), .QN(
        n36723) );
  DFF_X1 \DRAM_mem_reg[56][28]  ( .D(n7471), .CK(CLK), .Q(net253835), .QN(
        n36722) );
  DFF_X1 \DRAM_mem_reg[56][27]  ( .D(n7470), .CK(CLK), .Q(net253834), .QN(
        n36721) );
  DFF_X1 \DRAM_mem_reg[56][26]  ( .D(n7469), .CK(CLK), .Q(net253833), .QN(
        n36720) );
  DFF_X1 \DRAM_mem_reg[56][25]  ( .D(n7468), .CK(CLK), .Q(net253832), .QN(
        n36719) );
  DFF_X1 \DRAM_mem_reg[56][24]  ( .D(n7467), .CK(CLK), .Q(net253831), .QN(
        n36718) );
  DFF_X1 \DRAM_mem_reg[56][23]  ( .D(n7466), .CK(CLK), .Q(net253830), .QN(
        n36901) );
  DFF_X1 \DRAM_mem_reg[56][22]  ( .D(n7465), .CK(CLK), .Q(net253829), .QN(
        n36900) );
  DFF_X1 \DRAM_mem_reg[56][21]  ( .D(n7464), .CK(CLK), .Q(net253828), .QN(
        n36899) );
  DFF_X1 \DRAM_mem_reg[56][20]  ( .D(n7463), .CK(CLK), .Q(net253827), .QN(
        n36898) );
  DFF_X1 \DRAM_mem_reg[56][19]  ( .D(n7462), .CK(CLK), .Q(net253826), .QN(
        n36897) );
  DFF_X1 \DRAM_mem_reg[56][18]  ( .D(n7461), .CK(CLK), .Q(net253825), .QN(
        n36896) );
  DFF_X1 \DRAM_mem_reg[56][17]  ( .D(n7460), .CK(CLK), .Q(net253824), .QN(
        n36895) );
  DFF_X1 \DRAM_mem_reg[56][16]  ( .D(n7459), .CK(CLK), .Q(net253823), .QN(
        n36894) );
  DFF_X1 \DRAM_mem_reg[56][15]  ( .D(n7458), .CK(CLK), .Q(net253822), .QN(
        n36893) );
  DFF_X1 \DRAM_mem_reg[56][14]  ( .D(n7457), .CK(CLK), .Q(net253821), .QN(
        n36892) );
  DFF_X1 \DRAM_mem_reg[56][13]  ( .D(n7456), .CK(CLK), .Q(net253820), .QN(
        n36891) );
  DFF_X1 \DRAM_mem_reg[56][12]  ( .D(n7455), .CK(CLK), .Q(net253819), .QN(
        n36890) );
  DFF_X1 \DRAM_mem_reg[56][11]  ( .D(n7454), .CK(CLK), .Q(net253818), .QN(
        n36889) );
  DFF_X1 \DRAM_mem_reg[56][10]  ( .D(n7453), .CK(CLK), .Q(net253817), .QN(
        n36888) );
  DFF_X1 \DRAM_mem_reg[56][9]  ( .D(n7452), .CK(CLK), .Q(net253816), .QN(
        n36887) );
  DFF_X1 \DRAM_mem_reg[56][8]  ( .D(n7451), .CK(CLK), .Q(net253815), .QN(
        n36886) );
  DFF_X1 \DRAM_mem_reg[56][7]  ( .D(n7450), .CK(CLK), .Q(net253814), .QN(
        n36885) );
  DFF_X1 \DRAM_mem_reg[56][6]  ( .D(n7449), .CK(CLK), .Q(net253813), .QN(
        n36884) );
  DFF_X1 \DRAM_mem_reg[56][5]  ( .D(n7448), .CK(CLK), .Q(net253812), .QN(
        n36883) );
  DFF_X1 \DRAM_mem_reg[56][4]  ( .D(n7447), .CK(CLK), .Q(net253811), .QN(
        n36882) );
  DFF_X1 \DRAM_mem_reg[56][3]  ( .D(n7446), .CK(CLK), .Q(net253810), .QN(
        n36881) );
  DFF_X1 \DRAM_mem_reg[56][2]  ( .D(n7445), .CK(CLK), .Q(net253809), .QN(
        n36880) );
  DFF_X1 \DRAM_mem_reg[56][1]  ( .D(n7444), .CK(CLK), .Q(net253808), .QN(
        n36879) );
  DFF_X1 \DRAM_mem_reg[56][0]  ( .D(n7443), .CK(CLK), .Q(net253807), .QN(
        n36878) );
  DFF_X1 \DRAM_mem_reg[57][31]  ( .D(n7442), .CK(CLK), .QN(n35412) );
  DFF_X1 \DRAM_mem_reg[57][30]  ( .D(n7441), .CK(CLK), .QN(n35403) );
  DFF_X1 \DRAM_mem_reg[57][29]  ( .D(n7440), .CK(CLK), .QN(n35394) );
  DFF_X1 \DRAM_mem_reg[57][28]  ( .D(n7439), .CK(CLK), .QN(n35385) );
  DFF_X1 \DRAM_mem_reg[57][27]  ( .D(n7438), .CK(CLK), .QN(n35376) );
  DFF_X1 \DRAM_mem_reg[57][26]  ( .D(n7437), .CK(CLK), .QN(n35367) );
  DFF_X1 \DRAM_mem_reg[57][25]  ( .D(n7436), .CK(CLK), .QN(n35358) );
  DFF_X1 \DRAM_mem_reg[57][24]  ( .D(n7435), .CK(CLK), .QN(n35349) );
  DFF_X1 \DRAM_mem_reg[57][23]  ( .D(n7434), .CK(CLK), .QN(n35613) );
  DFF_X1 \DRAM_mem_reg[57][22]  ( .D(n7433), .CK(CLK), .QN(n35611) );
  DFF_X1 \DRAM_mem_reg[57][21]  ( .D(n7432), .CK(CLK), .QN(n35609) );
  DFF_X1 \DRAM_mem_reg[57][20]  ( .D(n7431), .CK(CLK), .QN(n35607) );
  DFF_X1 \DRAM_mem_reg[57][19]  ( .D(n7430), .CK(CLK), .QN(n35605) );
  DFF_X1 \DRAM_mem_reg[57][18]  ( .D(n7429), .CK(CLK), .QN(n35603) );
  DFF_X1 \DRAM_mem_reg[57][17]  ( .D(n7428), .CK(CLK), .QN(n35601) );
  DFF_X1 \DRAM_mem_reg[57][16]  ( .D(n7427), .CK(CLK), .QN(n35599) );
  DFF_X1 \DRAM_mem_reg[57][15]  ( .D(n7426), .CK(CLK), .QN(n35597) );
  DFF_X1 \DRAM_mem_reg[57][14]  ( .D(n7425), .CK(CLK), .QN(n35595) );
  DFF_X1 \DRAM_mem_reg[57][13]  ( .D(n7424), .CK(CLK), .QN(n35593) );
  DFF_X1 \DRAM_mem_reg[57][12]  ( .D(n7423), .CK(CLK), .QN(n35591) );
  DFF_X1 \DRAM_mem_reg[57][11]  ( .D(n7422), .CK(CLK), .QN(n35589) );
  DFF_X1 \DRAM_mem_reg[57][10]  ( .D(n7421), .CK(CLK), .QN(n35587) );
  DFF_X1 \DRAM_mem_reg[57][9]  ( .D(n7420), .CK(CLK), .QN(n35585) );
  DFF_X1 \DRAM_mem_reg[57][8]  ( .D(n7419), .CK(CLK), .QN(n35583) );
  DFF_X1 \DRAM_mem_reg[57][7]  ( .D(n7418), .CK(CLK), .QN(n35581) );
  DFF_X1 \DRAM_mem_reg[57][6]  ( .D(n7417), .CK(CLK), .QN(n35579) );
  DFF_X1 \DRAM_mem_reg[57][5]  ( .D(n7416), .CK(CLK), .QN(n35577) );
  DFF_X1 \DRAM_mem_reg[57][4]  ( .D(n7415), .CK(CLK), .QN(n35575) );
  DFF_X1 \DRAM_mem_reg[57][3]  ( .D(n7414), .CK(CLK), .QN(n35573) );
  DFF_X1 \DRAM_mem_reg[57][2]  ( .D(n7413), .CK(CLK), .QN(n35571) );
  DFF_X1 \DRAM_mem_reg[57][1]  ( .D(n7412), .CK(CLK), .QN(n35569) );
  DFF_X1 \DRAM_mem_reg[57][0]  ( .D(n7411), .CK(CLK), .QN(n35567) );
  DFF_X1 \DRAM_mem_reg[58][31]  ( .D(n7410), .CK(CLK), .QN(n35919) );
  DFF_X1 \DRAM_mem_reg[58][30]  ( .D(n7409), .CK(CLK), .QN(n35910) );
  DFF_X1 \DRAM_mem_reg[58][29]  ( .D(n7408), .CK(CLK), .QN(n35901) );
  DFF_X1 \DRAM_mem_reg[58][28]  ( .D(n7407), .CK(CLK), .QN(n35892) );
  DFF_X1 \DRAM_mem_reg[58][27]  ( .D(n7406), .CK(CLK), .QN(n35883) );
  DFF_X1 \DRAM_mem_reg[58][26]  ( .D(n7405), .CK(CLK), .QN(n35874) );
  DFF_X1 \DRAM_mem_reg[58][25]  ( .D(n7404), .CK(CLK), .QN(n35865) );
  DFF_X1 \DRAM_mem_reg[58][24]  ( .D(n7403), .CK(CLK), .QN(n35856) );
  DFF_X1 \DRAM_mem_reg[58][23]  ( .D(n7402), .CK(CLK), .QN(n36076) );
  DFF_X1 \DRAM_mem_reg[58][22]  ( .D(n7401), .CK(CLK), .QN(n36074) );
  DFF_X1 \DRAM_mem_reg[58][21]  ( .D(n7400), .CK(CLK), .QN(n36072) );
  DFF_X1 \DRAM_mem_reg[58][20]  ( .D(n7399), .CK(CLK), .QN(n36070) );
  DFF_X1 \DRAM_mem_reg[58][19]  ( .D(n7398), .CK(CLK), .QN(n36068) );
  DFF_X1 \DRAM_mem_reg[58][18]  ( .D(n7397), .CK(CLK), .QN(n36066) );
  DFF_X1 \DRAM_mem_reg[58][17]  ( .D(n7396), .CK(CLK), .QN(n36064) );
  DFF_X1 \DRAM_mem_reg[58][16]  ( .D(n7395), .CK(CLK), .QN(n36062) );
  DFF_X1 \DRAM_mem_reg[58][15]  ( .D(n7394), .CK(CLK), .QN(n36060) );
  DFF_X1 \DRAM_mem_reg[58][14]  ( .D(n7393), .CK(CLK), .QN(n36058) );
  DFF_X1 \DRAM_mem_reg[58][13]  ( .D(n7392), .CK(CLK), .QN(n36056) );
  DFF_X1 \DRAM_mem_reg[58][12]  ( .D(n7391), .CK(CLK), .QN(n36054) );
  DFF_X1 \DRAM_mem_reg[58][11]  ( .D(n7390), .CK(CLK), .QN(n36052) );
  DFF_X1 \DRAM_mem_reg[58][10]  ( .D(n7389), .CK(CLK), .QN(n36050) );
  DFF_X1 \DRAM_mem_reg[58][9]  ( .D(n7388), .CK(CLK), .QN(n36048) );
  DFF_X1 \DRAM_mem_reg[58][8]  ( .D(n7387), .CK(CLK), .QN(n36046) );
  DFF_X1 \DRAM_mem_reg[58][7]  ( .D(n7386), .CK(CLK), .QN(n36044) );
  DFF_X1 \DRAM_mem_reg[58][6]  ( .D(n7385), .CK(CLK), .QN(n36042) );
  DFF_X1 \DRAM_mem_reg[58][5]  ( .D(n7384), .CK(CLK), .QN(n36040) );
  DFF_X1 \DRAM_mem_reg[58][4]  ( .D(n7383), .CK(CLK), .QN(n36038) );
  DFF_X1 \DRAM_mem_reg[58][3]  ( .D(n7382), .CK(CLK), .QN(n36036) );
  DFF_X1 \DRAM_mem_reg[58][2]  ( .D(n7381), .CK(CLK), .QN(n36034) );
  DFF_X1 \DRAM_mem_reg[58][1]  ( .D(n7380), .CK(CLK), .QN(n36032) );
  DFF_X1 \DRAM_mem_reg[58][0]  ( .D(n7379), .CK(CLK), .QN(n36030) );
  DFF_X1 \DRAM_mem_reg[59][31]  ( .D(n7378), .CK(CLK), .Q(net253806), .QN(
        n37101) );
  DFF_X1 \DRAM_mem_reg[59][30]  ( .D(n7377), .CK(CLK), .Q(net253805), .QN(
        n37100) );
  DFF_X1 \DRAM_mem_reg[59][29]  ( .D(n7376), .CK(CLK), .Q(net253804), .QN(
        n37099) );
  DFF_X1 \DRAM_mem_reg[59][28]  ( .D(n7375), .CK(CLK), .Q(net253803), .QN(
        n37098) );
  DFF_X1 \DRAM_mem_reg[59][27]  ( .D(n7374), .CK(CLK), .Q(net253802), .QN(
        n37097) );
  DFF_X1 \DRAM_mem_reg[59][26]  ( .D(n7373), .CK(CLK), .Q(net253801), .QN(
        n37096) );
  DFF_X1 \DRAM_mem_reg[59][25]  ( .D(n7372), .CK(CLK), .Q(net253800), .QN(
        n37095) );
  DFF_X1 \DRAM_mem_reg[59][24]  ( .D(n7371), .CK(CLK), .Q(net253799), .QN(
        n37094) );
  DFF_X1 \DRAM_mem_reg[59][23]  ( .D(n7370), .CK(CLK), .Q(net253798), .QN(
        n37261) );
  DFF_X1 \DRAM_mem_reg[59][22]  ( .D(n7369), .CK(CLK), .Q(net253797), .QN(
        n37260) );
  DFF_X1 \DRAM_mem_reg[59][21]  ( .D(n7368), .CK(CLK), .Q(net253796), .QN(
        n37259) );
  DFF_X1 \DRAM_mem_reg[59][20]  ( .D(n7367), .CK(CLK), .Q(net253795), .QN(
        n37258) );
  DFF_X1 \DRAM_mem_reg[59][19]  ( .D(n7366), .CK(CLK), .Q(net253794), .QN(
        n37257) );
  DFF_X1 \DRAM_mem_reg[59][18]  ( .D(n7365), .CK(CLK), .Q(net253793), .QN(
        n37256) );
  DFF_X1 \DRAM_mem_reg[59][17]  ( .D(n7364), .CK(CLK), .Q(net253792), .QN(
        n37255) );
  DFF_X1 \DRAM_mem_reg[59][16]  ( .D(n7363), .CK(CLK), .Q(net253791), .QN(
        n37254) );
  DFF_X1 \DRAM_mem_reg[59][15]  ( .D(n7362), .CK(CLK), .Q(net253790), .QN(
        n37253) );
  DFF_X1 \DRAM_mem_reg[59][14]  ( .D(n7361), .CK(CLK), .Q(net253789), .QN(
        n37252) );
  DFF_X1 \DRAM_mem_reg[59][13]  ( .D(n7360), .CK(CLK), .Q(net253788), .QN(
        n37251) );
  DFF_X1 \DRAM_mem_reg[59][12]  ( .D(n7359), .CK(CLK), .Q(net253787), .QN(
        n37250) );
  DFF_X1 \DRAM_mem_reg[59][11]  ( .D(n7358), .CK(CLK), .Q(net253786), .QN(
        n37249) );
  DFF_X1 \DRAM_mem_reg[59][10]  ( .D(n7357), .CK(CLK), .Q(net253785), .QN(
        n37248) );
  DFF_X1 \DRAM_mem_reg[59][9]  ( .D(n7356), .CK(CLK), .Q(net253784), .QN(
        n37247) );
  DFF_X1 \DRAM_mem_reg[59][8]  ( .D(n7355), .CK(CLK), .Q(net253783), .QN(
        n37246) );
  DFF_X1 \DRAM_mem_reg[59][7]  ( .D(n7354), .CK(CLK), .Q(net253782), .QN(
        n37245) );
  DFF_X1 \DRAM_mem_reg[59][6]  ( .D(n7353), .CK(CLK), .Q(net253781), .QN(
        n37244) );
  DFF_X1 \DRAM_mem_reg[59][5]  ( .D(n7352), .CK(CLK), .Q(net253780), .QN(
        n37243) );
  DFF_X1 \DRAM_mem_reg[59][4]  ( .D(n7351), .CK(CLK), .Q(net253779), .QN(
        n37242) );
  DFF_X1 \DRAM_mem_reg[59][3]  ( .D(n7350), .CK(CLK), .Q(net253778), .QN(
        n37241) );
  DFF_X1 \DRAM_mem_reg[59][2]  ( .D(n7349), .CK(CLK), .Q(net253777), .QN(
        n37240) );
  DFF_X1 \DRAM_mem_reg[59][1]  ( .D(n7348), .CK(CLK), .Q(net253776), .QN(
        n37239) );
  DFF_X1 \DRAM_mem_reg[59][0]  ( .D(n7347), .CK(CLK), .Q(net253775), .QN(
        n37238) );
  DFF_X1 \DRAM_mem_reg[60][31]  ( .D(n7346), .CK(CLK), .QN(n36430) );
  DFF_X1 \DRAM_mem_reg[60][30]  ( .D(n7345), .CK(CLK), .QN(n36421) );
  DFF_X1 \DRAM_mem_reg[60][29]  ( .D(n7344), .CK(CLK), .QN(n36412) );
  DFF_X1 \DRAM_mem_reg[60][28]  ( .D(n7343), .CK(CLK), .QN(n36403) );
  DFF_X1 \DRAM_mem_reg[60][27]  ( .D(n7342), .CK(CLK), .QN(n36394) );
  DFF_X1 \DRAM_mem_reg[60][26]  ( .D(n7341), .CK(CLK), .QN(n36385) );
  DFF_X1 \DRAM_mem_reg[60][25]  ( .D(n7340), .CK(CLK), .QN(n36376) );
  DFF_X1 \DRAM_mem_reg[60][24]  ( .D(n7339), .CK(CLK), .QN(n36367) );
  DFF_X1 \DRAM_mem_reg[60][23]  ( .D(n7338), .CK(CLK), .QN(n36532) );
  DFF_X1 \DRAM_mem_reg[60][22]  ( .D(n7337), .CK(CLK), .QN(n36528) );
  DFF_X1 \DRAM_mem_reg[60][21]  ( .D(n7336), .CK(CLK), .QN(n36524) );
  DFF_X1 \DRAM_mem_reg[60][20]  ( .D(n7335), .CK(CLK), .QN(n36520) );
  DFF_X1 \DRAM_mem_reg[60][19]  ( .D(n7334), .CK(CLK), .QN(n36516) );
  DFF_X1 \DRAM_mem_reg[60][18]  ( .D(n7333), .CK(CLK), .QN(n36512) );
  DFF_X1 \DRAM_mem_reg[60][17]  ( .D(n7332), .CK(CLK), .QN(n36508) );
  DFF_X1 \DRAM_mem_reg[60][16]  ( .D(n7331), .CK(CLK), .QN(n36504) );
  DFF_X1 \DRAM_mem_reg[60][15]  ( .D(n7330), .CK(CLK), .QN(n36500) );
  DFF_X1 \DRAM_mem_reg[60][14]  ( .D(n7329), .CK(CLK), .QN(n36496) );
  DFF_X1 \DRAM_mem_reg[60][13]  ( .D(n7328), .CK(CLK), .QN(n36492) );
  DFF_X1 \DRAM_mem_reg[60][12]  ( .D(n7327), .CK(CLK), .QN(n36488) );
  DFF_X1 \DRAM_mem_reg[60][11]  ( .D(n7326), .CK(CLK), .QN(n36484) );
  DFF_X1 \DRAM_mem_reg[60][10]  ( .D(n7325), .CK(CLK), .QN(n36480) );
  DFF_X1 \DRAM_mem_reg[60][9]  ( .D(n7324), .CK(CLK), .QN(n36476) );
  DFF_X1 \DRAM_mem_reg[60][8]  ( .D(n7323), .CK(CLK), .QN(n36472) );
  DFF_X1 \DRAM_mem_reg[60][7]  ( .D(n7322), .CK(CLK), .QN(n36468) );
  DFF_X1 \DRAM_mem_reg[60][6]  ( .D(n7321), .CK(CLK), .QN(n36464) );
  DFF_X1 \DRAM_mem_reg[60][5]  ( .D(n7320), .CK(CLK), .QN(n36460) );
  DFF_X1 \DRAM_mem_reg[60][4]  ( .D(n7319), .CK(CLK), .QN(n36456) );
  DFF_X1 \DRAM_mem_reg[60][3]  ( .D(n7318), .CK(CLK), .QN(n36452) );
  DFF_X1 \DRAM_mem_reg[60][2]  ( .D(n7317), .CK(CLK), .QN(n36448) );
  DFF_X1 \DRAM_mem_reg[60][1]  ( .D(n7316), .CK(CLK), .QN(n36444) );
  DFF_X1 \DRAM_mem_reg[60][0]  ( .D(n7315), .CK(CLK), .QN(n36440) );
  DFF_X1 \DRAM_mem_reg[61][31]  ( .D(n7314), .CK(CLK), .Q(net253774), .QN(
        n36717) );
  DFF_X1 \DRAM_mem_reg[61][30]  ( .D(n7313), .CK(CLK), .Q(net253773), .QN(
        n36716) );
  DFF_X1 \DRAM_mem_reg[61][29]  ( .D(n7312), .CK(CLK), .Q(net253772), .QN(
        n36715) );
  DFF_X1 \DRAM_mem_reg[61][28]  ( .D(n7311), .CK(CLK), .Q(net253771), .QN(
        n36714) );
  DFF_X1 \DRAM_mem_reg[61][27]  ( .D(n7310), .CK(CLK), .Q(net253770), .QN(
        n36713) );
  DFF_X1 \DRAM_mem_reg[61][26]  ( .D(n7309), .CK(CLK), .Q(net253769), .QN(
        n36712) );
  DFF_X1 \DRAM_mem_reg[61][25]  ( .D(n7308), .CK(CLK), .Q(net253768), .QN(
        n36711) );
  DFF_X1 \DRAM_mem_reg[61][24]  ( .D(n7307), .CK(CLK), .Q(net253767), .QN(
        n36710) );
  DFF_X1 \DRAM_mem_reg[61][23]  ( .D(n7306), .CK(CLK), .Q(net253766), .QN(
        n36877) );
  DFF_X1 \DRAM_mem_reg[61][22]  ( .D(n7305), .CK(CLK), .Q(net253765), .QN(
        n36876) );
  DFF_X1 \DRAM_mem_reg[61][21]  ( .D(n7304), .CK(CLK), .Q(net253764), .QN(
        n36875) );
  DFF_X1 \DRAM_mem_reg[61][20]  ( .D(n7303), .CK(CLK), .Q(net253763), .QN(
        n36874) );
  DFF_X1 \DRAM_mem_reg[61][19]  ( .D(n7302), .CK(CLK), .Q(net253762), .QN(
        n36873) );
  DFF_X1 \DRAM_mem_reg[61][18]  ( .D(n7301), .CK(CLK), .Q(net253761), .QN(
        n36872) );
  DFF_X1 \DRAM_mem_reg[61][17]  ( .D(n7300), .CK(CLK), .Q(net253760), .QN(
        n36871) );
  DFF_X1 \DRAM_mem_reg[61][16]  ( .D(n7299), .CK(CLK), .Q(net253759), .QN(
        n36870) );
  DFF_X1 \DRAM_mem_reg[61][15]  ( .D(n7298), .CK(CLK), .Q(net253758), .QN(
        n36869) );
  DFF_X1 \DRAM_mem_reg[61][14]  ( .D(n7297), .CK(CLK), .Q(net253757), .QN(
        n36868) );
  DFF_X1 \DRAM_mem_reg[61][13]  ( .D(n7296), .CK(CLK), .Q(net253756), .QN(
        n36867) );
  DFF_X1 \DRAM_mem_reg[61][12]  ( .D(n7295), .CK(CLK), .Q(net253755), .QN(
        n36866) );
  DFF_X1 \DRAM_mem_reg[61][11]  ( .D(n7294), .CK(CLK), .Q(net253754), .QN(
        n36865) );
  DFF_X1 \DRAM_mem_reg[61][10]  ( .D(n7293), .CK(CLK), .Q(net253753), .QN(
        n36864) );
  DFF_X1 \DRAM_mem_reg[61][9]  ( .D(n7292), .CK(CLK), .Q(net253752), .QN(
        n36863) );
  DFF_X1 \DRAM_mem_reg[61][8]  ( .D(n7291), .CK(CLK), .Q(net253751), .QN(
        n36862) );
  DFF_X1 \DRAM_mem_reg[61][7]  ( .D(n7290), .CK(CLK), .Q(net253750), .QN(
        n36861) );
  DFF_X1 \DRAM_mem_reg[61][6]  ( .D(n7289), .CK(CLK), .Q(net253749), .QN(
        n36860) );
  DFF_X1 \DRAM_mem_reg[61][5]  ( .D(n7288), .CK(CLK), .Q(net253748), .QN(
        n36859) );
  DFF_X1 \DRAM_mem_reg[61][4]  ( .D(n7287), .CK(CLK), .Q(net253747), .QN(
        n36858) );
  DFF_X1 \DRAM_mem_reg[61][3]  ( .D(n7286), .CK(CLK), .Q(net253746), .QN(
        n36857) );
  DFF_X1 \DRAM_mem_reg[61][2]  ( .D(n7285), .CK(CLK), .Q(net253745), .QN(
        n36856) );
  DFF_X1 \DRAM_mem_reg[61][1]  ( .D(n7284), .CK(CLK), .Q(net253744), .QN(
        n36855) );
  DFF_X1 \DRAM_mem_reg[61][0]  ( .D(n7283), .CK(CLK), .Q(net253743), .QN(
        n36854) );
  DFF_X1 \DRAM_mem_reg[62][31]  ( .D(n7282), .CK(CLK), .QN(n35409) );
  DFF_X1 \DRAM_mem_reg[62][30]  ( .D(n7281), .CK(CLK), .QN(n35400) );
  DFF_X1 \DRAM_mem_reg[62][29]  ( .D(n7280), .CK(CLK), .QN(n35391) );
  DFF_X1 \DRAM_mem_reg[62][28]  ( .D(n7279), .CK(CLK), .QN(n35382) );
  DFF_X1 \DRAM_mem_reg[62][27]  ( .D(n7278), .CK(CLK), .QN(n35373) );
  DFF_X1 \DRAM_mem_reg[62][26]  ( .D(n7277), .CK(CLK), .QN(n35364) );
  DFF_X1 \DRAM_mem_reg[62][25]  ( .D(n7276), .CK(CLK), .QN(n35355) );
  DFF_X1 \DRAM_mem_reg[62][24]  ( .D(n7275), .CK(CLK), .QN(n35346) );
  DFF_X1 \DRAM_mem_reg[62][23]  ( .D(n7274), .CK(CLK), .QN(n35660) );
  DFF_X1 \DRAM_mem_reg[62][22]  ( .D(n7273), .CK(CLK), .QN(n35658) );
  DFF_X1 \DRAM_mem_reg[62][21]  ( .D(n7272), .CK(CLK), .QN(n35656) );
  DFF_X1 \DRAM_mem_reg[62][20]  ( .D(n7271), .CK(CLK), .QN(n35654) );
  DFF_X1 \DRAM_mem_reg[62][19]  ( .D(n7270), .CK(CLK), .QN(n35652) );
  DFF_X1 \DRAM_mem_reg[62][18]  ( .D(n7269), .CK(CLK), .QN(n35650) );
  DFF_X1 \DRAM_mem_reg[62][17]  ( .D(n7268), .CK(CLK), .QN(n35648) );
  DFF_X1 \DRAM_mem_reg[62][16]  ( .D(n7267), .CK(CLK), .QN(n35646) );
  DFF_X1 \DRAM_mem_reg[62][15]  ( .D(n7266), .CK(CLK), .QN(n35644) );
  DFF_X1 \DRAM_mem_reg[62][14]  ( .D(n7265), .CK(CLK), .QN(n35642) );
  DFF_X1 \DRAM_mem_reg[62][13]  ( .D(n7264), .CK(CLK), .QN(n35640) );
  DFF_X1 \DRAM_mem_reg[62][12]  ( .D(n7263), .CK(CLK), .QN(n35638) );
  DFF_X1 \DRAM_mem_reg[62][11]  ( .D(n7262), .CK(CLK), .QN(n35636) );
  DFF_X1 \DRAM_mem_reg[62][10]  ( .D(n7261), .CK(CLK), .QN(n35634) );
  DFF_X1 \DRAM_mem_reg[62][9]  ( .D(n7260), .CK(CLK), .QN(n35632) );
  DFF_X1 \DRAM_mem_reg[62][8]  ( .D(n7259), .CK(CLK), .QN(n35630) );
  DFF_X1 \DRAM_mem_reg[62][7]  ( .D(n7258), .CK(CLK), .QN(n35628) );
  DFF_X1 \DRAM_mem_reg[62][6]  ( .D(n7257), .CK(CLK), .QN(n35626) );
  DFF_X1 \DRAM_mem_reg[62][5]  ( .D(n7256), .CK(CLK), .QN(n35624) );
  DFF_X1 \DRAM_mem_reg[62][4]  ( .D(n7255), .CK(CLK), .QN(n35622) );
  DFF_X1 \DRAM_mem_reg[62][3]  ( .D(n7254), .CK(CLK), .QN(n35620) );
  DFF_X1 \DRAM_mem_reg[62][2]  ( .D(n7253), .CK(CLK), .QN(n35618) );
  DFF_X1 \DRAM_mem_reg[62][1]  ( .D(n7252), .CK(CLK), .QN(n35616) );
  DFF_X1 \DRAM_mem_reg[62][0]  ( .D(n7251), .CK(CLK), .QN(n35614) );
  DFF_X1 \DRAM_mem_reg[63][31]  ( .D(n7250), .CK(CLK), .QN(n35920) );
  DFF_X1 \DRAM_mem_reg[63][30]  ( .D(n7249), .CK(CLK), .QN(n35911) );
  DFF_X1 \DRAM_mem_reg[63][29]  ( .D(n7248), .CK(CLK), .QN(n35902) );
  DFF_X1 \DRAM_mem_reg[63][28]  ( .D(n7247), .CK(CLK), .QN(n35893) );
  DFF_X1 \DRAM_mem_reg[63][27]  ( .D(n7246), .CK(CLK), .QN(n35884) );
  DFF_X1 \DRAM_mem_reg[63][26]  ( .D(n7245), .CK(CLK), .QN(n35875) );
  DFF_X1 \DRAM_mem_reg[63][25]  ( .D(n7244), .CK(CLK), .QN(n35866) );
  DFF_X1 \DRAM_mem_reg[63][24]  ( .D(n7243), .CK(CLK), .QN(n35857) );
  DFF_X1 \DRAM_mem_reg[63][23]  ( .D(n7242), .CK(CLK), .QN(n36124) );
  DFF_X1 \DRAM_mem_reg[63][22]  ( .D(n7241), .CK(CLK), .QN(n36122) );
  DFF_X1 \DRAM_mem_reg[63][21]  ( .D(n7240), .CK(CLK), .QN(n36120) );
  DFF_X1 \DRAM_mem_reg[63][20]  ( .D(n7239), .CK(CLK), .QN(n36118) );
  DFF_X1 \DRAM_mem_reg[63][19]  ( .D(n7238), .CK(CLK), .QN(n36116) );
  DFF_X1 \DRAM_mem_reg[63][18]  ( .D(n7237), .CK(CLK), .QN(n36114) );
  DFF_X1 \DRAM_mem_reg[63][17]  ( .D(n7236), .CK(CLK), .QN(n36112) );
  DFF_X1 \DRAM_mem_reg[63][16]  ( .D(n7235), .CK(CLK), .QN(n36110) );
  DFF_X1 \DRAM_mem_reg[63][15]  ( .D(n7234), .CK(CLK), .QN(n36108) );
  DFF_X1 \DRAM_mem_reg[63][14]  ( .D(n7233), .CK(CLK), .QN(n36106) );
  DFF_X1 \DRAM_mem_reg[63][13]  ( .D(n7232), .CK(CLK), .QN(n36104) );
  DFF_X1 \DRAM_mem_reg[63][12]  ( .D(n7231), .CK(CLK), .QN(n36102) );
  DFF_X1 \DRAM_mem_reg[63][11]  ( .D(n7230), .CK(CLK), .QN(n36100) );
  DFF_X1 \DRAM_mem_reg[63][10]  ( .D(n7229), .CK(CLK), .QN(n36098) );
  DFF_X1 \DRAM_mem_reg[63][9]  ( .D(n7228), .CK(CLK), .QN(n36096) );
  DFF_X1 \DRAM_mem_reg[63][8]  ( .D(n7227), .CK(CLK), .QN(n36094) );
  DFF_X1 \DRAM_mem_reg[63][7]  ( .D(n7226), .CK(CLK), .QN(n36092) );
  DFF_X1 \DRAM_mem_reg[63][6]  ( .D(n7225), .CK(CLK), .QN(n36090) );
  DFF_X1 \DRAM_mem_reg[63][5]  ( .D(n7224), .CK(CLK), .QN(n36088) );
  DFF_X1 \DRAM_mem_reg[63][4]  ( .D(n7223), .CK(CLK), .QN(n36086) );
  DFF_X1 \DRAM_mem_reg[63][3]  ( .D(n7222), .CK(CLK), .QN(n36084) );
  DFF_X1 \DRAM_mem_reg[63][2]  ( .D(n7221), .CK(CLK), .QN(n36082) );
  DFF_X1 \DRAM_mem_reg[63][1]  ( .D(n7220), .CK(CLK), .QN(n36080) );
  DFF_X1 \DRAM_mem_reg[63][0]  ( .D(n7219), .CK(CLK), .QN(n36078) );
  DFF_X1 \DRAM_mem_reg[64][31]  ( .D(n7218), .CK(CLK), .Q(n5558), .QN(n36709)
         );
  DFF_X1 \DRAM_mem_reg[64][30]  ( .D(n7217), .CK(CLK), .Q(n5608), .QN(n36708)
         );
  DFF_X1 \DRAM_mem_reg[64][29]  ( .D(n7216), .CK(CLK), .Q(n5650), .QN(n36707)
         );
  DFF_X1 \DRAM_mem_reg[64][28]  ( .D(n7215), .CK(CLK), .Q(n5692), .QN(n36706)
         );
  DFF_X1 \DRAM_mem_reg[64][27]  ( .D(n7214), .CK(CLK), .Q(n5734), .QN(n36705)
         );
  DFF_X1 \DRAM_mem_reg[64][26]  ( .D(n7213), .CK(CLK), .Q(n5776), .QN(n36704)
         );
  DFF_X1 \DRAM_mem_reg[64][25]  ( .D(n7212), .CK(CLK), .Q(n5818), .QN(n36703)
         );
  DFF_X1 \DRAM_mem_reg[64][24]  ( .D(n7211), .CK(CLK), .Q(n5860), .QN(n36702)
         );
  DFF_X1 \DRAM_mem_reg[64][23]  ( .D(n7210), .CK(CLK), .Q(n5902), .QN(n36853)
         );
  DFF_X1 \DRAM_mem_reg[64][22]  ( .D(n7209), .CK(CLK), .Q(n5944), .QN(n36852)
         );
  DFF_X1 \DRAM_mem_reg[64][21]  ( .D(n7208), .CK(CLK), .Q(n5986), .QN(n36851)
         );
  DFF_X1 \DRAM_mem_reg[64][20]  ( .D(n7207), .CK(CLK), .Q(n6028), .QN(n36850)
         );
  DFF_X1 \DRAM_mem_reg[64][19]  ( .D(n7206), .CK(CLK), .Q(n6070), .QN(n36849)
         );
  DFF_X1 \DRAM_mem_reg[64][18]  ( .D(n7205), .CK(CLK), .Q(n6112), .QN(n36848)
         );
  DFF_X1 \DRAM_mem_reg[64][17]  ( .D(n7204), .CK(CLK), .Q(n6154), .QN(n36847)
         );
  DFF_X1 \DRAM_mem_reg[64][16]  ( .D(n7203), .CK(CLK), .Q(n6196), .QN(n36846)
         );
  DFF_X1 \DRAM_mem_reg[64][15]  ( .D(n7202), .CK(CLK), .Q(n6238), .QN(n36845)
         );
  DFF_X1 \DRAM_mem_reg[64][14]  ( .D(n7201), .CK(CLK), .Q(n6280), .QN(n36844)
         );
  DFF_X1 \DRAM_mem_reg[64][13]  ( .D(n7200), .CK(CLK), .Q(n6322), .QN(n36843)
         );
  DFF_X1 \DRAM_mem_reg[64][12]  ( .D(n7199), .CK(CLK), .Q(n6364), .QN(n36842)
         );
  DFF_X1 \DRAM_mem_reg[64][11]  ( .D(n7198), .CK(CLK), .Q(n6534), .QN(n36841)
         );
  DFF_X1 \DRAM_mem_reg[64][10]  ( .D(n7197), .CK(CLK), .Q(n6576), .QN(n36840)
         );
  DFF_X1 \DRAM_mem_reg[64][9]  ( .D(n7196), .CK(CLK), .Q(n6618), .QN(n36839)
         );
  DFF_X1 \DRAM_mem_reg[64][8]  ( .D(n7195), .CK(CLK), .Q(n6660), .QN(n36838)
         );
  DFF_X1 \DRAM_mem_reg[64][7]  ( .D(n7194), .CK(CLK), .Q(n9294), .QN(n36837)
         );
  DFF_X1 \DRAM_mem_reg[64][6]  ( .D(n7193), .CK(CLK), .Q(n9336), .QN(n36836)
         );
  DFF_X1 \DRAM_mem_reg[64][5]  ( .D(n7192), .CK(CLK), .Q(n9378), .QN(n36835)
         );
  DFF_X1 \DRAM_mem_reg[64][4]  ( .D(n7191), .CK(CLK), .Q(n9420), .QN(n36834)
         );
  DFF_X1 \DRAM_mem_reg[64][3]  ( .D(n7190), .CK(CLK), .Q(n9462), .QN(n36833)
         );
  DFF_X1 \DRAM_mem_reg[64][2]  ( .D(n7189), .CK(CLK), .Q(n9504), .QN(n36832)
         );
  DFF_X1 \DRAM_mem_reg[64][1]  ( .D(n7188), .CK(CLK), .Q(n9546), .QN(n36831)
         );
  DFF_X1 \DRAM_mem_reg[64][0]  ( .D(n7187), .CK(CLK), .Q(n9609), .QN(n36830)
         );
  DFF_X1 \DRAM_mem_reg[65][31]  ( .D(n7186), .CK(CLK), .QN(n35677) );
  DFF_X1 \DRAM_mem_reg[65][30]  ( .D(n7185), .CK(CLK), .QN(n35676) );
  DFF_X1 \DRAM_mem_reg[65][29]  ( .D(n7184), .CK(CLK), .QN(n35675) );
  DFF_X1 \DRAM_mem_reg[65][28]  ( .D(n7183), .CK(CLK), .QN(n35674) );
  DFF_X1 \DRAM_mem_reg[65][27]  ( .D(n7182), .CK(CLK), .QN(n35673) );
  DFF_X1 \DRAM_mem_reg[65][26]  ( .D(n7181), .CK(CLK), .QN(n35672) );
  DFF_X1 \DRAM_mem_reg[65][25]  ( .D(n7180), .CK(CLK), .QN(n35671) );
  DFF_X1 \DRAM_mem_reg[65][24]  ( .D(n7179), .CK(CLK), .QN(n35670) );
  DFF_X1 \DRAM_mem_reg[65][23]  ( .D(n7178), .CK(CLK), .QN(n35757) );
  DFF_X1 \DRAM_mem_reg[65][22]  ( .D(n7177), .CK(CLK), .QN(n35756) );
  DFF_X1 \DRAM_mem_reg[65][21]  ( .D(n7176), .CK(CLK), .QN(n35755) );
  DFF_X1 \DRAM_mem_reg[65][20]  ( .D(n7175), .CK(CLK), .QN(n35754) );
  DFF_X1 \DRAM_mem_reg[65][19]  ( .D(n7174), .CK(CLK), .QN(n35753) );
  DFF_X1 \DRAM_mem_reg[65][18]  ( .D(n7173), .CK(CLK), .QN(n35752) );
  DFF_X1 \DRAM_mem_reg[65][17]  ( .D(n7172), .CK(CLK), .QN(n35751) );
  DFF_X1 \DRAM_mem_reg[65][16]  ( .D(n7171), .CK(CLK), .QN(n35750) );
  DFF_X1 \DRAM_mem_reg[65][15]  ( .D(n7170), .CK(CLK), .QN(n35749) );
  DFF_X1 \DRAM_mem_reg[65][14]  ( .D(n7169), .CK(CLK), .QN(n35748) );
  DFF_X1 \DRAM_mem_reg[65][13]  ( .D(n7168), .CK(CLK), .QN(n35747) );
  DFF_X1 \DRAM_mem_reg[65][12]  ( .D(n7167), .CK(CLK), .QN(n35746) );
  DFF_X1 \DRAM_mem_reg[65][11]  ( .D(n7166), .CK(CLK), .QN(n35745) );
  DFF_X1 \DRAM_mem_reg[65][10]  ( .D(n7165), .CK(CLK), .QN(n35744) );
  DFF_X1 \DRAM_mem_reg[65][9]  ( .D(n7164), .CK(CLK), .QN(n35743) );
  DFF_X1 \DRAM_mem_reg[65][8]  ( .D(n7163), .CK(CLK), .QN(n35742) );
  DFF_X1 \DRAM_mem_reg[65][7]  ( .D(n7162), .CK(CLK), .QN(n35741) );
  DFF_X1 \DRAM_mem_reg[65][6]  ( .D(n7161), .CK(CLK), .QN(n35740) );
  DFF_X1 \DRAM_mem_reg[65][5]  ( .D(n7160), .CK(CLK), .QN(n35739) );
  DFF_X1 \DRAM_mem_reg[65][4]  ( .D(n7159), .CK(CLK), .QN(n35738) );
  DFF_X1 \DRAM_mem_reg[65][3]  ( .D(n7158), .CK(CLK), .QN(n35737) );
  DFF_X1 \DRAM_mem_reg[65][2]  ( .D(n7157), .CK(CLK), .QN(n35736) );
  DFF_X1 \DRAM_mem_reg[65][1]  ( .D(n7156), .CK(CLK), .QN(n35735) );
  DFF_X1 \DRAM_mem_reg[65][0]  ( .D(n7155), .CK(CLK), .QN(n35734) );
  DFF_X1 \DRAM_mem_reg[66][31]  ( .D(n7154), .CK(CLK), .QN(n36189) );
  DFF_X1 \DRAM_mem_reg[66][30]  ( .D(n7153), .CK(CLK), .QN(n36188) );
  DFF_X1 \DRAM_mem_reg[66][29]  ( .D(n7152), .CK(CLK), .QN(n36187) );
  DFF_X1 \DRAM_mem_reg[66][28]  ( .D(n7151), .CK(CLK), .QN(n36186) );
  DFF_X1 \DRAM_mem_reg[66][27]  ( .D(n7150), .CK(CLK), .QN(n36185) );
  DFF_X1 \DRAM_mem_reg[66][26]  ( .D(n7149), .CK(CLK), .QN(n36184) );
  DFF_X1 \DRAM_mem_reg[66][25]  ( .D(n7148), .CK(CLK), .QN(n36183) );
  DFF_X1 \DRAM_mem_reg[66][24]  ( .D(n7147), .CK(CLK), .QN(n36182) );
  DFF_X1 \DRAM_mem_reg[66][23]  ( .D(n7146), .CK(CLK), .QN(n36269) );
  DFF_X1 \DRAM_mem_reg[66][22]  ( .D(n7145), .CK(CLK), .QN(n36268) );
  DFF_X1 \DRAM_mem_reg[66][21]  ( .D(n7144), .CK(CLK), .QN(n36267) );
  DFF_X1 \DRAM_mem_reg[66][20]  ( .D(n7143), .CK(CLK), .QN(n36266) );
  DFF_X1 \DRAM_mem_reg[66][19]  ( .D(n7142), .CK(CLK), .QN(n36265) );
  DFF_X1 \DRAM_mem_reg[66][18]  ( .D(n7141), .CK(CLK), .QN(n36264) );
  DFF_X1 \DRAM_mem_reg[66][17]  ( .D(n7140), .CK(CLK), .QN(n36263) );
  DFF_X1 \DRAM_mem_reg[66][16]  ( .D(n7139), .CK(CLK), .QN(n36262) );
  DFF_X1 \DRAM_mem_reg[66][15]  ( .D(n7138), .CK(CLK), .QN(n36261) );
  DFF_X1 \DRAM_mem_reg[66][14]  ( .D(n7137), .CK(CLK), .QN(n36260) );
  DFF_X1 \DRAM_mem_reg[66][13]  ( .D(n7136), .CK(CLK), .QN(n36259) );
  DFF_X1 \DRAM_mem_reg[66][12]  ( .D(n7135), .CK(CLK), .QN(n36258) );
  DFF_X1 \DRAM_mem_reg[66][11]  ( .D(n7134), .CK(CLK), .QN(n36257) );
  DFF_X1 \DRAM_mem_reg[66][10]  ( .D(n7133), .CK(CLK), .QN(n36256) );
  DFF_X1 \DRAM_mem_reg[66][9]  ( .D(n7132), .CK(CLK), .QN(n36255) );
  DFF_X1 \DRAM_mem_reg[66][8]  ( .D(n7131), .CK(CLK), .QN(n36254) );
  DFF_X1 \DRAM_mem_reg[66][7]  ( .D(n7130), .CK(CLK), .QN(n36253) );
  DFF_X1 \DRAM_mem_reg[66][6]  ( .D(n7129), .CK(CLK), .QN(n36252) );
  DFF_X1 \DRAM_mem_reg[66][5]  ( .D(n7128), .CK(CLK), .QN(n36251) );
  DFF_X1 \DRAM_mem_reg[66][4]  ( .D(n7127), .CK(CLK), .QN(n36250) );
  DFF_X1 \DRAM_mem_reg[66][3]  ( .D(n7126), .CK(CLK), .QN(n36249) );
  DFF_X1 \DRAM_mem_reg[66][2]  ( .D(n7125), .CK(CLK), .QN(n36248) );
  DFF_X1 \DRAM_mem_reg[66][1]  ( .D(n7124), .CK(CLK), .QN(n36247) );
  DFF_X1 \DRAM_mem_reg[66][0]  ( .D(n7123), .CK(CLK), .QN(n36246) );
  DFF_X1 \DRAM_mem_reg[67][31]  ( .D(n7122), .CK(CLK), .QN(n35165) );
  DFF_X1 \DRAM_mem_reg[67][30]  ( .D(n7121), .CK(CLK), .QN(n35164) );
  DFF_X1 \DRAM_mem_reg[67][29]  ( .D(n7120), .CK(CLK), .QN(n35163) );
  DFF_X1 \DRAM_mem_reg[67][28]  ( .D(n7119), .CK(CLK), .QN(n35162) );
  DFF_X1 \DRAM_mem_reg[67][27]  ( .D(n7118), .CK(CLK), .QN(n35161) );
  DFF_X1 \DRAM_mem_reg[67][26]  ( .D(n7117), .CK(CLK), .QN(n35160) );
  DFF_X1 \DRAM_mem_reg[67][25]  ( .D(n7116), .CK(CLK), .QN(n35159) );
  DFF_X1 \DRAM_mem_reg[67][24]  ( .D(n7115), .CK(CLK), .QN(n35158) );
  DFF_X1 \DRAM_mem_reg[67][23]  ( .D(n7114), .CK(CLK), .QN(n35245) );
  DFF_X1 \DRAM_mem_reg[67][22]  ( .D(n7113), .CK(CLK), .QN(n35244) );
  DFF_X1 \DRAM_mem_reg[67][21]  ( .D(n7112), .CK(CLK), .QN(n35243) );
  DFF_X1 \DRAM_mem_reg[67][20]  ( .D(n7111), .CK(CLK), .QN(n35242) );
  DFF_X1 \DRAM_mem_reg[67][19]  ( .D(n7110), .CK(CLK), .QN(n35241) );
  DFF_X1 \DRAM_mem_reg[67][18]  ( .D(n7109), .CK(CLK), .QN(n35240) );
  DFF_X1 \DRAM_mem_reg[67][17]  ( .D(n7108), .CK(CLK), .QN(n35239) );
  DFF_X1 \DRAM_mem_reg[67][16]  ( .D(n7107), .CK(CLK), .QN(n35238) );
  DFF_X1 \DRAM_mem_reg[67][15]  ( .D(n7106), .CK(CLK), .QN(n35237) );
  DFF_X1 \DRAM_mem_reg[67][14]  ( .D(n7105), .CK(CLK), .QN(n35236) );
  DFF_X1 \DRAM_mem_reg[67][13]  ( .D(n7104), .CK(CLK), .QN(n35235) );
  DFF_X1 \DRAM_mem_reg[67][12]  ( .D(n7103), .CK(CLK), .QN(n35234) );
  DFF_X1 \DRAM_mem_reg[67][11]  ( .D(n7102), .CK(CLK), .QN(n35233) );
  DFF_X1 \DRAM_mem_reg[67][10]  ( .D(n7101), .CK(CLK), .QN(n35232) );
  DFF_X1 \DRAM_mem_reg[67][9]  ( .D(n7100), .CK(CLK), .QN(n35231) );
  DFF_X1 \DRAM_mem_reg[67][8]  ( .D(n7099), .CK(CLK), .QN(n35230) );
  DFF_X1 \DRAM_mem_reg[67][7]  ( .D(n7098), .CK(CLK), .QN(n35229) );
  DFF_X1 \DRAM_mem_reg[67][6]  ( .D(n7097), .CK(CLK), .QN(n35228) );
  DFF_X1 \DRAM_mem_reg[67][5]  ( .D(n7096), .CK(CLK), .QN(n35227) );
  DFF_X1 \DRAM_mem_reg[67][4]  ( .D(n7095), .CK(CLK), .QN(n35226) );
  DFF_X1 \DRAM_mem_reg[67][3]  ( .D(n7094), .CK(CLK), .QN(n35225) );
  DFF_X1 \DRAM_mem_reg[67][2]  ( .D(n7093), .CK(CLK), .QN(n35224) );
  DFF_X1 \DRAM_mem_reg[67][1]  ( .D(n7092), .CK(CLK), .QN(n35223) );
  DFF_X1 \DRAM_mem_reg[67][0]  ( .D(n7091), .CK(CLK), .QN(n35222) );
  DFF_X1 \DRAM_mem_reg[68][31]  ( .D(n7090), .CK(CLK), .Q(net253742), .QN(
        n37093) );
  DFF_X1 \DRAM_mem_reg[68][30]  ( .D(n7089), .CK(CLK), .Q(net253741), .QN(
        n37092) );
  DFF_X1 \DRAM_mem_reg[68][29]  ( .D(n7088), .CK(CLK), .Q(net253740), .QN(
        n37091) );
  DFF_X1 \DRAM_mem_reg[68][28]  ( .D(n7087), .CK(CLK), .Q(net253739), .QN(
        n37090) );
  DFF_X1 \DRAM_mem_reg[68][27]  ( .D(n7086), .CK(CLK), .Q(net253738), .QN(
        n37089) );
  DFF_X1 \DRAM_mem_reg[68][26]  ( .D(n7085), .CK(CLK), .Q(net253737), .QN(
        n37088) );
  DFF_X1 \DRAM_mem_reg[68][25]  ( .D(n7084), .CK(CLK), .Q(net253736), .QN(
        n37087) );
  DFF_X1 \DRAM_mem_reg[68][24]  ( .D(n7083), .CK(CLK), .Q(net253735), .QN(
        n37086) );
  DFF_X1 \DRAM_mem_reg[68][23]  ( .D(n7082), .CK(CLK), .Q(net253734), .QN(
        n37237) );
  DFF_X1 \DRAM_mem_reg[68][22]  ( .D(n7081), .CK(CLK), .Q(net253733), .QN(
        n37236) );
  DFF_X1 \DRAM_mem_reg[68][21]  ( .D(n7080), .CK(CLK), .Q(net253732), .QN(
        n37235) );
  DFF_X1 \DRAM_mem_reg[68][20]  ( .D(n7079), .CK(CLK), .Q(net253731), .QN(
        n37234) );
  DFF_X1 \DRAM_mem_reg[68][19]  ( .D(n7078), .CK(CLK), .Q(net253730), .QN(
        n37233) );
  DFF_X1 \DRAM_mem_reg[68][18]  ( .D(n7077), .CK(CLK), .Q(net253729), .QN(
        n37232) );
  DFF_X1 \DRAM_mem_reg[68][17]  ( .D(n7076), .CK(CLK), .Q(net253728), .QN(
        n37231) );
  DFF_X1 \DRAM_mem_reg[68][16]  ( .D(n7075), .CK(CLK), .Q(net253727), .QN(
        n37230) );
  DFF_X1 \DRAM_mem_reg[68][15]  ( .D(n7074), .CK(CLK), .Q(net253726), .QN(
        n37229) );
  DFF_X1 \DRAM_mem_reg[68][14]  ( .D(n7073), .CK(CLK), .Q(net253725), .QN(
        n37228) );
  DFF_X1 \DRAM_mem_reg[68][13]  ( .D(n7072), .CK(CLK), .Q(net253724), .QN(
        n37227) );
  DFF_X1 \DRAM_mem_reg[68][12]  ( .D(n7071), .CK(CLK), .Q(net253723), .QN(
        n37226) );
  DFF_X1 \DRAM_mem_reg[68][11]  ( .D(n7070), .CK(CLK), .Q(net253722), .QN(
        n37225) );
  DFF_X1 \DRAM_mem_reg[68][10]  ( .D(n7069), .CK(CLK), .Q(net253721), .QN(
        n37224) );
  DFF_X1 \DRAM_mem_reg[68][9]  ( .D(n7068), .CK(CLK), .Q(net253720), .QN(
        n37223) );
  DFF_X1 \DRAM_mem_reg[68][8]  ( .D(n7067), .CK(CLK), .Q(net253719), .QN(
        n37222) );
  DFF_X1 \DRAM_mem_reg[68][7]  ( .D(n7066), .CK(CLK), .Q(net253718), .QN(
        n37221) );
  DFF_X1 \DRAM_mem_reg[68][6]  ( .D(n7065), .CK(CLK), .Q(net253717), .QN(
        n37220) );
  DFF_X1 \DRAM_mem_reg[68][5]  ( .D(n7064), .CK(CLK), .Q(net253716), .QN(
        n37219) );
  DFF_X1 \DRAM_mem_reg[68][4]  ( .D(n7063), .CK(CLK), .Q(net253715), .QN(
        n37218) );
  DFF_X1 \DRAM_mem_reg[68][3]  ( .D(n7062), .CK(CLK), .Q(net253714), .QN(
        n37217) );
  DFF_X1 \DRAM_mem_reg[68][2]  ( .D(n7061), .CK(CLK), .Q(net253713), .QN(
        n37216) );
  DFF_X1 \DRAM_mem_reg[68][1]  ( .D(n7060), .CK(CLK), .Q(net253712), .QN(
        n37215) );
  DFF_X1 \DRAM_mem_reg[68][0]  ( .D(n7059), .CK(CLK), .Q(net253711), .QN(
        n37214) );
  DFF_X1 \DRAM_mem_reg[69][31]  ( .D(n7058), .CK(CLK), .Q(net253710), .QN(
        n36701) );
  DFF_X1 \DRAM_mem_reg[69][30]  ( .D(n7057), .CK(CLK), .Q(net253709), .QN(
        n36700) );
  DFF_X1 \DRAM_mem_reg[69][29]  ( .D(n7056), .CK(CLK), .Q(net253708), .QN(
        n36699) );
  DFF_X1 \DRAM_mem_reg[69][28]  ( .D(n7055), .CK(CLK), .Q(net253707), .QN(
        n36698) );
  DFF_X1 \DRAM_mem_reg[69][27]  ( .D(n7054), .CK(CLK), .Q(net253706), .QN(
        n36697) );
  DFF_X1 \DRAM_mem_reg[69][26]  ( .D(n7053), .CK(CLK), .Q(net253705), .QN(
        n36696) );
  DFF_X1 \DRAM_mem_reg[69][25]  ( .D(n7052), .CK(CLK), .Q(net253704), .QN(
        n36695) );
  DFF_X1 \DRAM_mem_reg[69][24]  ( .D(n7051), .CK(CLK), .Q(net253703), .QN(
        n36694) );
  DFF_X1 \DRAM_mem_reg[69][23]  ( .D(n7050), .CK(CLK), .Q(net253702), .QN(
        n36829) );
  DFF_X1 \DRAM_mem_reg[69][22]  ( .D(n7049), .CK(CLK), .Q(net253701), .QN(
        n36828) );
  DFF_X1 \DRAM_mem_reg[69][21]  ( .D(n7048), .CK(CLK), .Q(net253700), .QN(
        n36827) );
  DFF_X1 \DRAM_mem_reg[69][20]  ( .D(n7047), .CK(CLK), .Q(net253699), .QN(
        n36826) );
  DFF_X1 \DRAM_mem_reg[69][19]  ( .D(n7046), .CK(CLK), .Q(net253698), .QN(
        n36825) );
  DFF_X1 \DRAM_mem_reg[69][18]  ( .D(n7045), .CK(CLK), .Q(net253697), .QN(
        n36824) );
  DFF_X1 \DRAM_mem_reg[69][17]  ( .D(n7044), .CK(CLK), .Q(net253696), .QN(
        n36823) );
  DFF_X1 \DRAM_mem_reg[69][16]  ( .D(n7043), .CK(CLK), .Q(net253695), .QN(
        n36822) );
  DFF_X1 \DRAM_mem_reg[69][15]  ( .D(n7042), .CK(CLK), .Q(net253694), .QN(
        n36821) );
  DFF_X1 \DRAM_mem_reg[69][14]  ( .D(n7041), .CK(CLK), .Q(net253693), .QN(
        n36820) );
  DFF_X1 \DRAM_mem_reg[69][13]  ( .D(n7040), .CK(CLK), .Q(net253692), .QN(
        n36819) );
  DFF_X1 \DRAM_mem_reg[69][12]  ( .D(n7039), .CK(CLK), .Q(net253691), .QN(
        n36818) );
  DFF_X1 \DRAM_mem_reg[69][11]  ( .D(n7038), .CK(CLK), .Q(net253690), .QN(
        n36817) );
  DFF_X1 \DRAM_mem_reg[69][10]  ( .D(n7037), .CK(CLK), .Q(net253689), .QN(
        n36816) );
  DFF_X1 \DRAM_mem_reg[69][9]  ( .D(n7036), .CK(CLK), .Q(net253688), .QN(
        n36815) );
  DFF_X1 \DRAM_mem_reg[69][8]  ( .D(n7035), .CK(CLK), .Q(net253687), .QN(
        n36814) );
  DFF_X1 \DRAM_mem_reg[69][7]  ( .D(n7034), .CK(CLK), .Q(net253686), .QN(
        n36813) );
  DFF_X1 \DRAM_mem_reg[69][6]  ( .D(n7033), .CK(CLK), .Q(net253685), .QN(
        n36812) );
  DFF_X1 \DRAM_mem_reg[69][5]  ( .D(n7032), .CK(CLK), .Q(net253684), .QN(
        n36811) );
  DFF_X1 \DRAM_mem_reg[69][4]  ( .D(n7031), .CK(CLK), .Q(net253683), .QN(
        n36810) );
  DFF_X1 \DRAM_mem_reg[69][3]  ( .D(n7030), .CK(CLK), .Q(net253682), .QN(
        n36809) );
  DFF_X1 \DRAM_mem_reg[69][2]  ( .D(n7029), .CK(CLK), .Q(net253681), .QN(
        n36808) );
  DFF_X1 \DRAM_mem_reg[69][1]  ( .D(n7028), .CK(CLK), .Q(net253680), .QN(
        n36807) );
  DFF_X1 \DRAM_mem_reg[69][0]  ( .D(n7027), .CK(CLK), .Q(net253679), .QN(
        n36806) );
  DFF_X1 \DRAM_mem_reg[70][31]  ( .D(n7026), .CK(CLK), .QN(n35669) );
  DFF_X1 \DRAM_mem_reg[70][30]  ( .D(n7025), .CK(CLK), .QN(n35668) );
  DFF_X1 \DRAM_mem_reg[70][29]  ( .D(n7024), .CK(CLK), .QN(n35667) );
  DFF_X1 \DRAM_mem_reg[70][28]  ( .D(n7023), .CK(CLK), .QN(n35666) );
  DFF_X1 \DRAM_mem_reg[70][27]  ( .D(n7022), .CK(CLK), .QN(n35665) );
  DFF_X1 \DRAM_mem_reg[70][26]  ( .D(n7021), .CK(CLK), .QN(n35664) );
  DFF_X1 \DRAM_mem_reg[70][25]  ( .D(n7020), .CK(CLK), .QN(n35663) );
  DFF_X1 \DRAM_mem_reg[70][24]  ( .D(n7019), .CK(CLK), .QN(n35662) );
  DFF_X1 \DRAM_mem_reg[70][23]  ( .D(n7018), .CK(CLK), .QN(n35733) );
  DFF_X1 \DRAM_mem_reg[70][22]  ( .D(n7017), .CK(CLK), .QN(n35732) );
  DFF_X1 \DRAM_mem_reg[70][21]  ( .D(n7016), .CK(CLK), .QN(n35731) );
  DFF_X1 \DRAM_mem_reg[70][20]  ( .D(n7015), .CK(CLK), .QN(n35730) );
  DFF_X1 \DRAM_mem_reg[70][19]  ( .D(n7014), .CK(CLK), .QN(n35729) );
  DFF_X1 \DRAM_mem_reg[70][18]  ( .D(n7013), .CK(CLK), .QN(n35728) );
  DFF_X1 \DRAM_mem_reg[70][17]  ( .D(n7012), .CK(CLK), .QN(n35727) );
  DFF_X1 \DRAM_mem_reg[70][16]  ( .D(n7011), .CK(CLK), .QN(n35726) );
  DFF_X1 \DRAM_mem_reg[70][15]  ( .D(n7010), .CK(CLK), .QN(n35725) );
  DFF_X1 \DRAM_mem_reg[70][14]  ( .D(n7009), .CK(CLK), .QN(n35724) );
  DFF_X1 \DRAM_mem_reg[70][13]  ( .D(n7008), .CK(CLK), .QN(n35723) );
  DFF_X1 \DRAM_mem_reg[70][12]  ( .D(n7007), .CK(CLK), .QN(n35722) );
  DFF_X1 \DRAM_mem_reg[70][11]  ( .D(n7006), .CK(CLK), .QN(n35721) );
  DFF_X1 \DRAM_mem_reg[70][10]  ( .D(n7005), .CK(CLK), .QN(n35720) );
  DFF_X1 \DRAM_mem_reg[70][9]  ( .D(n7004), .CK(CLK), .QN(n35719) );
  DFF_X1 \DRAM_mem_reg[70][8]  ( .D(n7003), .CK(CLK), .QN(n35718) );
  DFF_X1 \DRAM_mem_reg[70][7]  ( .D(n7002), .CK(CLK), .QN(n35717) );
  DFF_X1 \DRAM_mem_reg[70][6]  ( .D(n7001), .CK(CLK), .QN(n35716) );
  DFF_X1 \DRAM_mem_reg[70][5]  ( .D(n7000), .CK(CLK), .QN(n35715) );
  DFF_X1 \DRAM_mem_reg[70][4]  ( .D(n6999), .CK(CLK), .QN(n35714) );
  DFF_X1 \DRAM_mem_reg[70][3]  ( .D(n6998), .CK(CLK), .QN(n35713) );
  DFF_X1 \DRAM_mem_reg[70][2]  ( .D(n6997), .CK(CLK), .QN(n35712) );
  DFF_X1 \DRAM_mem_reg[70][1]  ( .D(n6996), .CK(CLK), .QN(n35711) );
  DFF_X1 \DRAM_mem_reg[70][0]  ( .D(n6995), .CK(CLK), .QN(n35710) );
  DFF_X1 \DRAM_mem_reg[71][31]  ( .D(n6994), .CK(CLK), .QN(n36181) );
  DFF_X1 \DRAM_mem_reg[71][30]  ( .D(n6993), .CK(CLK), .QN(n36180) );
  DFF_X1 \DRAM_mem_reg[71][29]  ( .D(n6992), .CK(CLK), .QN(n36179) );
  DFF_X1 \DRAM_mem_reg[71][28]  ( .D(n6991), .CK(CLK), .QN(n36178) );
  DFF_X1 \DRAM_mem_reg[71][27]  ( .D(n6990), .CK(CLK), .QN(n36177) );
  DFF_X1 \DRAM_mem_reg[71][26]  ( .D(n6989), .CK(CLK), .QN(n36176) );
  DFF_X1 \DRAM_mem_reg[71][25]  ( .D(n6988), .CK(CLK), .QN(n36175) );
  DFF_X1 \DRAM_mem_reg[71][24]  ( .D(n6987), .CK(CLK), .QN(n36174) );
  DFF_X1 \DRAM_mem_reg[71][23]  ( .D(n6986), .CK(CLK), .QN(n36245) );
  DFF_X1 \DRAM_mem_reg[71][22]  ( .D(n6985), .CK(CLK), .QN(n36244) );
  DFF_X1 \DRAM_mem_reg[71][21]  ( .D(n6984), .CK(CLK), .QN(n36243) );
  DFF_X1 \DRAM_mem_reg[71][20]  ( .D(n6983), .CK(CLK), .QN(n36242) );
  DFF_X1 \DRAM_mem_reg[71][19]  ( .D(n6982), .CK(CLK), .QN(n36241) );
  DFF_X1 \DRAM_mem_reg[71][18]  ( .D(n6981), .CK(CLK), .QN(n36240) );
  DFF_X1 \DRAM_mem_reg[71][17]  ( .D(n6980), .CK(CLK), .QN(n36239) );
  DFF_X1 \DRAM_mem_reg[71][16]  ( .D(n6979), .CK(CLK), .QN(n36238) );
  DFF_X1 \DRAM_mem_reg[71][15]  ( .D(n6978), .CK(CLK), .QN(n36237) );
  DFF_X1 \DRAM_mem_reg[71][14]  ( .D(n6977), .CK(CLK), .QN(n36236) );
  DFF_X1 \DRAM_mem_reg[71][13]  ( .D(n6976), .CK(CLK), .QN(n36235) );
  DFF_X1 \DRAM_mem_reg[71][12]  ( .D(n6975), .CK(CLK), .QN(n36234) );
  DFF_X1 \DRAM_mem_reg[71][11]  ( .D(n6974), .CK(CLK), .QN(n36233) );
  DFF_X1 \DRAM_mem_reg[71][10]  ( .D(n6973), .CK(CLK), .QN(n36232) );
  DFF_X1 \DRAM_mem_reg[71][9]  ( .D(n6972), .CK(CLK), .QN(n36231) );
  DFF_X1 \DRAM_mem_reg[71][8]  ( .D(n6971), .CK(CLK), .QN(n36230) );
  DFF_X1 \DRAM_mem_reg[71][7]  ( .D(n6970), .CK(CLK), .QN(n36229) );
  DFF_X1 \DRAM_mem_reg[71][6]  ( .D(n6969), .CK(CLK), .QN(n36228) );
  DFF_X1 \DRAM_mem_reg[71][5]  ( .D(n6968), .CK(CLK), .QN(n36227) );
  DFF_X1 \DRAM_mem_reg[71][4]  ( .D(n6967), .CK(CLK), .QN(n36226) );
  DFF_X1 \DRAM_mem_reg[71][3]  ( .D(n6966), .CK(CLK), .QN(n36225) );
  DFF_X1 \DRAM_mem_reg[71][2]  ( .D(n6965), .CK(CLK), .QN(n36224) );
  DFF_X1 \DRAM_mem_reg[71][1]  ( .D(n6964), .CK(CLK), .QN(n36223) );
  DFF_X1 \DRAM_mem_reg[71][0]  ( .D(n6963), .CK(CLK), .QN(n36222) );
  DFF_X1 \DRAM_mem_reg[72][31]  ( .D(n6962), .CK(CLK), .QN(n35157) );
  DFF_X1 \DRAM_mem_reg[72][30]  ( .D(n6961), .CK(CLK), .QN(n35156) );
  DFF_X1 \DRAM_mem_reg[72][29]  ( .D(n6960), .CK(CLK), .QN(n35155) );
  DFF_X1 \DRAM_mem_reg[72][28]  ( .D(n6959), .CK(CLK), .QN(n35154) );
  DFF_X1 \DRAM_mem_reg[72][27]  ( .D(n6958), .CK(CLK), .QN(n35153) );
  DFF_X1 \DRAM_mem_reg[72][26]  ( .D(n6957), .CK(CLK), .QN(n35152) );
  DFF_X1 \DRAM_mem_reg[72][25]  ( .D(n6956), .CK(CLK), .QN(n35151) );
  DFF_X1 \DRAM_mem_reg[72][24]  ( .D(n6955), .CK(CLK), .QN(n35150) );
  DFF_X1 \DRAM_mem_reg[72][23]  ( .D(n6954), .CK(CLK), .QN(n35221) );
  DFF_X1 \DRAM_mem_reg[72][22]  ( .D(n6953), .CK(CLK), .QN(n35220) );
  DFF_X1 \DRAM_mem_reg[72][21]  ( .D(n6952), .CK(CLK), .QN(n35219) );
  DFF_X1 \DRAM_mem_reg[72][20]  ( .D(n6951), .CK(CLK), .QN(n35218) );
  DFF_X1 \DRAM_mem_reg[72][19]  ( .D(n6950), .CK(CLK), .QN(n35217) );
  DFF_X1 \DRAM_mem_reg[72][18]  ( .D(n6949), .CK(CLK), .QN(n35216) );
  DFF_X1 \DRAM_mem_reg[72][17]  ( .D(n6948), .CK(CLK), .QN(n35215) );
  DFF_X1 \DRAM_mem_reg[72][16]  ( .D(n6947), .CK(CLK), .QN(n35214) );
  DFF_X1 \DRAM_mem_reg[72][15]  ( .D(n6946), .CK(CLK), .QN(n35213) );
  DFF_X1 \DRAM_mem_reg[72][14]  ( .D(n6945), .CK(CLK), .QN(n35212) );
  DFF_X1 \DRAM_mem_reg[72][13]  ( .D(n6944), .CK(CLK), .QN(n35211) );
  DFF_X1 \DRAM_mem_reg[72][12]  ( .D(n6943), .CK(CLK), .QN(n35210) );
  DFF_X1 \DRAM_mem_reg[72][11]  ( .D(n6942), .CK(CLK), .QN(n35209) );
  DFF_X1 \DRAM_mem_reg[72][10]  ( .D(n6941), .CK(CLK), .QN(n35208) );
  DFF_X1 \DRAM_mem_reg[72][9]  ( .D(n6940), .CK(CLK), .QN(n35207) );
  DFF_X1 \DRAM_mem_reg[72][8]  ( .D(n6939), .CK(CLK), .QN(n35206) );
  DFF_X1 \DRAM_mem_reg[72][7]  ( .D(n6938), .CK(CLK), .QN(n35205) );
  DFF_X1 \DRAM_mem_reg[72][6]  ( .D(n6937), .CK(CLK), .QN(n35204) );
  DFF_X1 \DRAM_mem_reg[72][5]  ( .D(n6936), .CK(CLK), .QN(n35203) );
  DFF_X1 \DRAM_mem_reg[72][4]  ( .D(n6935), .CK(CLK), .QN(n35202) );
  DFF_X1 \DRAM_mem_reg[72][3]  ( .D(n6934), .CK(CLK), .QN(n35201) );
  DFF_X1 \DRAM_mem_reg[72][2]  ( .D(n6933), .CK(CLK), .QN(n35200) );
  DFF_X1 \DRAM_mem_reg[72][1]  ( .D(n6932), .CK(CLK), .QN(n35199) );
  DFF_X1 \DRAM_mem_reg[72][0]  ( .D(n6931), .CK(CLK), .QN(n35198) );
  DFF_X1 \DRAM_mem_reg[73][31]  ( .D(n6930), .CK(CLK), .Q(net253678), .QN(
        n37085) );
  DFF_X1 \DRAM_mem_reg[73][30]  ( .D(n6929), .CK(CLK), .Q(net253677), .QN(
        n37084) );
  DFF_X1 \DRAM_mem_reg[73][29]  ( .D(n6928), .CK(CLK), .Q(net253676), .QN(
        n37083) );
  DFF_X1 \DRAM_mem_reg[73][28]  ( .D(n6927), .CK(CLK), .Q(net253675), .QN(
        n37082) );
  DFF_X1 \DRAM_mem_reg[73][27]  ( .D(n6926), .CK(CLK), .Q(net253674), .QN(
        n37081) );
  DFF_X1 \DRAM_mem_reg[73][26]  ( .D(n6925), .CK(CLK), .Q(net253673), .QN(
        n37080) );
  DFF_X1 \DRAM_mem_reg[73][25]  ( .D(n6924), .CK(CLK), .Q(net253672), .QN(
        n37079) );
  DFF_X1 \DRAM_mem_reg[73][24]  ( .D(n6923), .CK(CLK), .Q(net253671), .QN(
        n37078) );
  DFF_X1 \DRAM_mem_reg[73][23]  ( .D(n6922), .CK(CLK), .Q(net253670), .QN(
        n37213) );
  DFF_X1 \DRAM_mem_reg[73][22]  ( .D(n6921), .CK(CLK), .Q(net253669), .QN(
        n37212) );
  DFF_X1 \DRAM_mem_reg[73][21]  ( .D(n6920), .CK(CLK), .Q(net253668), .QN(
        n37211) );
  DFF_X1 \DRAM_mem_reg[73][20]  ( .D(n6919), .CK(CLK), .Q(net253667), .QN(
        n37210) );
  DFF_X1 \DRAM_mem_reg[73][19]  ( .D(n6918), .CK(CLK), .Q(net253666), .QN(
        n37209) );
  DFF_X1 \DRAM_mem_reg[73][18]  ( .D(n6917), .CK(CLK), .Q(net253665), .QN(
        n37208) );
  DFF_X1 \DRAM_mem_reg[73][17]  ( .D(n6916), .CK(CLK), .Q(net253664), .QN(
        n37207) );
  DFF_X1 \DRAM_mem_reg[73][16]  ( .D(n6915), .CK(CLK), .Q(net253663), .QN(
        n37206) );
  DFF_X1 \DRAM_mem_reg[73][15]  ( .D(n6914), .CK(CLK), .Q(net253662), .QN(
        n37205) );
  DFF_X1 \DRAM_mem_reg[73][14]  ( .D(n6913), .CK(CLK), .Q(net253661), .QN(
        n37204) );
  DFF_X1 \DRAM_mem_reg[73][13]  ( .D(n6912), .CK(CLK), .Q(net253660), .QN(
        n37203) );
  DFF_X1 \DRAM_mem_reg[73][12]  ( .D(n6911), .CK(CLK), .Q(net253659), .QN(
        n37202) );
  DFF_X1 \DRAM_mem_reg[73][11]  ( .D(n6910), .CK(CLK), .Q(net253658), .QN(
        n37201) );
  DFF_X1 \DRAM_mem_reg[73][10]  ( .D(n6909), .CK(CLK), .Q(net253657), .QN(
        n37200) );
  DFF_X1 \DRAM_mem_reg[73][9]  ( .D(n6908), .CK(CLK), .Q(net253656), .QN(
        n37199) );
  DFF_X1 \DRAM_mem_reg[73][8]  ( .D(n6907), .CK(CLK), .Q(net253655), .QN(
        n37198) );
  DFF_X1 \DRAM_mem_reg[73][7]  ( .D(n6906), .CK(CLK), .Q(net253654), .QN(
        n37197) );
  DFF_X1 \DRAM_mem_reg[73][6]  ( .D(n6905), .CK(CLK), .Q(net253653), .QN(
        n37196) );
  DFF_X1 \DRAM_mem_reg[73][5]  ( .D(n6904), .CK(CLK), .Q(net253652), .QN(
        n37195) );
  DFF_X1 \DRAM_mem_reg[73][4]  ( .D(n6903), .CK(CLK), .Q(net253651), .QN(
        n37194) );
  DFF_X1 \DRAM_mem_reg[73][3]  ( .D(n6902), .CK(CLK), .Q(net253650), .QN(
        n37193) );
  DFF_X1 \DRAM_mem_reg[73][2]  ( .D(n6901), .CK(CLK), .Q(net253649), .QN(
        n37192) );
  DFF_X1 \DRAM_mem_reg[73][1]  ( .D(n6900), .CK(CLK), .Q(net253648), .QN(
        n37191) );
  DFF_X1 \DRAM_mem_reg[73][0]  ( .D(n6899), .CK(CLK), .Q(net253647), .QN(
        n37190) );
  DFF_X1 \DRAM_mem_reg[74][31]  ( .D(n6898), .CK(CLK), .Q(net253646), .QN(
        n36693) );
  DFF_X1 \DRAM_mem_reg[74][30]  ( .D(n6897), .CK(CLK), .Q(net253645), .QN(
        n36692) );
  DFF_X1 \DRAM_mem_reg[74][29]  ( .D(n6896), .CK(CLK), .Q(net253644), .QN(
        n36691) );
  DFF_X1 \DRAM_mem_reg[74][28]  ( .D(n6895), .CK(CLK), .Q(net253643), .QN(
        n36690) );
  DFF_X1 \DRAM_mem_reg[74][27]  ( .D(n6894), .CK(CLK), .Q(net253642), .QN(
        n36689) );
  DFF_X1 \DRAM_mem_reg[74][26]  ( .D(n6893), .CK(CLK), .Q(net253641), .QN(
        n36688) );
  DFF_X1 \DRAM_mem_reg[74][25]  ( .D(n6892), .CK(CLK), .Q(net253640), .QN(
        n36687) );
  DFF_X1 \DRAM_mem_reg[74][24]  ( .D(n6891), .CK(CLK), .Q(net253639), .QN(
        n36686) );
  DFF_X1 \DRAM_mem_reg[74][23]  ( .D(n6890), .CK(CLK), .Q(net253638), .QN(
        n36805) );
  DFF_X1 \DRAM_mem_reg[74][22]  ( .D(n6889), .CK(CLK), .Q(net253637), .QN(
        n36804) );
  DFF_X1 \DRAM_mem_reg[74][21]  ( .D(n6888), .CK(CLK), .Q(net253636), .QN(
        n36803) );
  DFF_X1 \DRAM_mem_reg[74][20]  ( .D(n6887), .CK(CLK), .Q(net253635), .QN(
        n36802) );
  DFF_X1 \DRAM_mem_reg[74][19]  ( .D(n6886), .CK(CLK), .Q(net253634), .QN(
        n36801) );
  DFF_X1 \DRAM_mem_reg[74][18]  ( .D(n6885), .CK(CLK), .Q(net253633), .QN(
        n36800) );
  DFF_X1 \DRAM_mem_reg[74][17]  ( .D(n6884), .CK(CLK), .Q(net253632), .QN(
        n36799) );
  DFF_X1 \DRAM_mem_reg[74][16]  ( .D(n6883), .CK(CLK), .Q(net253631), .QN(
        n36798) );
  DFF_X1 \DRAM_mem_reg[74][15]  ( .D(n6882), .CK(CLK), .Q(net253630), .QN(
        n36797) );
  DFF_X1 \DRAM_mem_reg[74][14]  ( .D(n6881), .CK(CLK), .Q(net253629), .QN(
        n36796) );
  DFF_X1 \DRAM_mem_reg[74][13]  ( .D(n6880), .CK(CLK), .Q(net253628), .QN(
        n36795) );
  DFF_X1 \DRAM_mem_reg[74][12]  ( .D(n6879), .CK(CLK), .Q(net253627), .QN(
        n36794) );
  DFF_X1 \DRAM_mem_reg[74][11]  ( .D(n6878), .CK(CLK), .Q(net253626), .QN(
        n36793) );
  DFF_X1 \DRAM_mem_reg[74][10]  ( .D(n6877), .CK(CLK), .Q(net253625), .QN(
        n36792) );
  DFF_X1 \DRAM_mem_reg[74][9]  ( .D(n6876), .CK(CLK), .Q(net253624), .QN(
        n36791) );
  DFF_X1 \DRAM_mem_reg[74][8]  ( .D(n6875), .CK(CLK), .Q(net253623), .QN(
        n36790) );
  DFF_X1 \DRAM_mem_reg[74][7]  ( .D(n6874), .CK(CLK), .Q(net253622), .QN(
        n36789) );
  DFF_X1 \DRAM_mem_reg[74][6]  ( .D(n6873), .CK(CLK), .Q(net253621), .QN(
        n36788) );
  DFF_X1 \DRAM_mem_reg[74][5]  ( .D(n6872), .CK(CLK), .Q(net253620), .QN(
        n36787) );
  DFF_X1 \DRAM_mem_reg[74][4]  ( .D(n6871), .CK(CLK), .Q(net253619), .QN(
        n36786) );
  DFF_X1 \DRAM_mem_reg[74][3]  ( .D(n6870), .CK(CLK), .Q(net253618), .QN(
        n36785) );
  DFF_X1 \DRAM_mem_reg[74][2]  ( .D(n6869), .CK(CLK), .Q(net253617), .QN(
        n36784) );
  DFF_X1 \DRAM_mem_reg[74][1]  ( .D(n6868), .CK(CLK), .Q(net253616), .QN(
        n36783) );
  DFF_X1 \DRAM_mem_reg[74][0]  ( .D(n6867), .CK(CLK), .Q(net253615), .QN(
        n36782) );
  DFF_X1 \DRAM_mem_reg[75][31]  ( .D(n6866), .CK(CLK), .QN(n35917) );
  DFF_X1 \DRAM_mem_reg[75][30]  ( .D(n6865), .CK(CLK), .QN(n35908) );
  DFF_X1 \DRAM_mem_reg[75][29]  ( .D(n6864), .CK(CLK), .QN(n35899) );
  DFF_X1 \DRAM_mem_reg[75][28]  ( .D(n6863), .CK(CLK), .QN(n35890) );
  DFF_X1 \DRAM_mem_reg[75][27]  ( .D(n6862), .CK(CLK), .QN(n35881) );
  DFF_X1 \DRAM_mem_reg[75][26]  ( .D(n6861), .CK(CLK), .QN(n35872) );
  DFF_X1 \DRAM_mem_reg[75][25]  ( .D(n6860), .CK(CLK), .QN(n35863) );
  DFF_X1 \DRAM_mem_reg[75][24]  ( .D(n6859), .CK(CLK), .QN(n35854) );
  DFF_X1 \DRAM_mem_reg[75][23]  ( .D(n6858), .CK(CLK), .QN(n36018) );
  DFF_X1 \DRAM_mem_reg[75][22]  ( .D(n6857), .CK(CLK), .QN(n36014) );
  DFF_X1 \DRAM_mem_reg[75][21]  ( .D(n6856), .CK(CLK), .QN(n36010) );
  DFF_X1 \DRAM_mem_reg[75][20]  ( .D(n6855), .CK(CLK), .QN(n36006) );
  DFF_X1 \DRAM_mem_reg[75][19]  ( .D(n6854), .CK(CLK), .QN(n36002) );
  DFF_X1 \DRAM_mem_reg[75][18]  ( .D(n6853), .CK(CLK), .QN(n35998) );
  DFF_X1 \DRAM_mem_reg[75][17]  ( .D(n6852), .CK(CLK), .QN(n35994) );
  DFF_X1 \DRAM_mem_reg[75][16]  ( .D(n6851), .CK(CLK), .QN(n35990) );
  DFF_X1 \DRAM_mem_reg[75][15]  ( .D(n6850), .CK(CLK), .QN(n35986) );
  DFF_X1 \DRAM_mem_reg[75][14]  ( .D(n6849), .CK(CLK), .QN(n35982) );
  DFF_X1 \DRAM_mem_reg[75][13]  ( .D(n6848), .CK(CLK), .QN(n35978) );
  DFF_X1 \DRAM_mem_reg[75][12]  ( .D(n6847), .CK(CLK), .QN(n35974) );
  DFF_X1 \DRAM_mem_reg[75][11]  ( .D(n6846), .CK(CLK), .QN(n35970) );
  DFF_X1 \DRAM_mem_reg[75][10]  ( .D(n6845), .CK(CLK), .QN(n35966) );
  DFF_X1 \DRAM_mem_reg[75][9]  ( .D(n6844), .CK(CLK), .QN(n35962) );
  DFF_X1 \DRAM_mem_reg[75][8]  ( .D(n6843), .CK(CLK), .QN(n35958) );
  DFF_X1 \DRAM_mem_reg[75][7]  ( .D(n6842), .CK(CLK), .QN(n35954) );
  DFF_X1 \DRAM_mem_reg[75][6]  ( .D(n6841), .CK(CLK), .QN(n35950) );
  DFF_X1 \DRAM_mem_reg[75][5]  ( .D(n6840), .CK(CLK), .QN(n35946) );
  DFF_X1 \DRAM_mem_reg[75][4]  ( .D(n6839), .CK(CLK), .QN(n35942) );
  DFF_X1 \DRAM_mem_reg[75][3]  ( .D(n6838), .CK(CLK), .QN(n35938) );
  DFF_X1 \DRAM_mem_reg[75][2]  ( .D(n6837), .CK(CLK), .QN(n35934) );
  DFF_X1 \DRAM_mem_reg[75][1]  ( .D(n6836), .CK(CLK), .QN(n35930) );
  DFF_X1 \DRAM_mem_reg[75][0]  ( .D(n6835), .CK(CLK), .QN(n35926) );
  DFF_X1 \DRAM_mem_reg[76][31]  ( .D(n6834), .CK(CLK), .QN(n36429) );
  DFF_X1 \DRAM_mem_reg[76][30]  ( .D(n6833), .CK(CLK), .QN(n36420) );
  DFF_X1 \DRAM_mem_reg[76][29]  ( .D(n6832), .CK(CLK), .QN(n36411) );
  DFF_X1 \DRAM_mem_reg[76][28]  ( .D(n6831), .CK(CLK), .QN(n36402) );
  DFF_X1 \DRAM_mem_reg[76][27]  ( .D(n6830), .CK(CLK), .QN(n36393) );
  DFF_X1 \DRAM_mem_reg[76][26]  ( .D(n6829), .CK(CLK), .QN(n36384) );
  DFF_X1 \DRAM_mem_reg[76][25]  ( .D(n6828), .CK(CLK), .QN(n36375) );
  DFF_X1 \DRAM_mem_reg[76][24]  ( .D(n6827), .CK(CLK), .QN(n36366) );
  DFF_X1 \DRAM_mem_reg[76][23]  ( .D(n6826), .CK(CLK), .QN(n36530) );
  DFF_X1 \DRAM_mem_reg[76][22]  ( .D(n6825), .CK(CLK), .QN(n36526) );
  DFF_X1 \DRAM_mem_reg[76][21]  ( .D(n6824), .CK(CLK), .QN(n36522) );
  DFF_X1 \DRAM_mem_reg[76][20]  ( .D(n6823), .CK(CLK), .QN(n36518) );
  DFF_X1 \DRAM_mem_reg[76][19]  ( .D(n6822), .CK(CLK), .QN(n36514) );
  DFF_X1 \DRAM_mem_reg[76][18]  ( .D(n6821), .CK(CLK), .QN(n36510) );
  DFF_X1 \DRAM_mem_reg[76][17]  ( .D(n6820), .CK(CLK), .QN(n36506) );
  DFF_X1 \DRAM_mem_reg[76][16]  ( .D(n6819), .CK(CLK), .QN(n36502) );
  DFF_X1 \DRAM_mem_reg[76][15]  ( .D(n6818), .CK(CLK), .QN(n36498) );
  DFF_X1 \DRAM_mem_reg[76][14]  ( .D(n6817), .CK(CLK), .QN(n36494) );
  DFF_X1 \DRAM_mem_reg[76][13]  ( .D(n6816), .CK(CLK), .QN(n36490) );
  DFF_X1 \DRAM_mem_reg[76][12]  ( .D(n6815), .CK(CLK), .QN(n36486) );
  DFF_X1 \DRAM_mem_reg[76][11]  ( .D(n6814), .CK(CLK), .QN(n36482) );
  DFF_X1 \DRAM_mem_reg[76][10]  ( .D(n6813), .CK(CLK), .QN(n36478) );
  DFF_X1 \DRAM_mem_reg[76][9]  ( .D(n6812), .CK(CLK), .QN(n36474) );
  DFF_X1 \DRAM_mem_reg[76][8]  ( .D(n6811), .CK(CLK), .QN(n36470) );
  DFF_X1 \DRAM_mem_reg[76][7]  ( .D(n6810), .CK(CLK), .QN(n36466) );
  DFF_X1 \DRAM_mem_reg[76][6]  ( .D(n6809), .CK(CLK), .QN(n36462) );
  DFF_X1 \DRAM_mem_reg[76][5]  ( .D(n6808), .CK(CLK), .QN(n36458) );
  DFF_X1 \DRAM_mem_reg[76][4]  ( .D(n6807), .CK(CLK), .QN(n36454) );
  DFF_X1 \DRAM_mem_reg[76][3]  ( .D(n6806), .CK(CLK), .QN(n36450) );
  DFF_X1 \DRAM_mem_reg[76][2]  ( .D(n6805), .CK(CLK), .QN(n36446) );
  DFF_X1 \DRAM_mem_reg[76][1]  ( .D(n6804), .CK(CLK), .QN(n36442) );
  DFF_X1 \DRAM_mem_reg[76][0]  ( .D(n6803), .CK(CLK), .QN(n36438) );
  DFF_X1 \DRAM_mem_reg[77][31]  ( .D(n6802), .CK(CLK), .QN(n35405) );
  DFF_X1 \DRAM_mem_reg[77][30]  ( .D(n6801), .CK(CLK), .QN(n35396) );
  DFF_X1 \DRAM_mem_reg[77][29]  ( .D(n6800), .CK(CLK), .QN(n35387) );
  DFF_X1 \DRAM_mem_reg[77][28]  ( .D(n6799), .CK(CLK), .QN(n35378) );
  DFF_X1 \DRAM_mem_reg[77][27]  ( .D(n6798), .CK(CLK), .QN(n35369) );
  DFF_X1 \DRAM_mem_reg[77][26]  ( .D(n6797), .CK(CLK), .QN(n35360) );
  DFF_X1 \DRAM_mem_reg[77][25]  ( .D(n6796), .CK(CLK), .QN(n35351) );
  DFF_X1 \DRAM_mem_reg[77][24]  ( .D(n6795), .CK(CLK), .QN(n35342) );
  DFF_X1 \DRAM_mem_reg[77][23]  ( .D(n6794), .CK(CLK), .QN(n35506) );
  DFF_X1 \DRAM_mem_reg[77][22]  ( .D(n6793), .CK(CLK), .QN(n35502) );
  DFF_X1 \DRAM_mem_reg[77][21]  ( .D(n6792), .CK(CLK), .QN(n35498) );
  DFF_X1 \DRAM_mem_reg[77][20]  ( .D(n6791), .CK(CLK), .QN(n35494) );
  DFF_X1 \DRAM_mem_reg[77][19]  ( .D(n6790), .CK(CLK), .QN(n35490) );
  DFF_X1 \DRAM_mem_reg[77][18]  ( .D(n6789), .CK(CLK), .QN(n35486) );
  DFF_X1 \DRAM_mem_reg[77][17]  ( .D(n6788), .CK(CLK), .QN(n35482) );
  DFF_X1 \DRAM_mem_reg[77][16]  ( .D(n6787), .CK(CLK), .QN(n35478) );
  DFF_X1 \DRAM_mem_reg[77][15]  ( .D(n6786), .CK(CLK), .QN(n35474) );
  DFF_X1 \DRAM_mem_reg[77][14]  ( .D(n6785), .CK(CLK), .QN(n35470) );
  DFF_X1 \DRAM_mem_reg[77][13]  ( .D(n6784), .CK(CLK), .QN(n35466) );
  DFF_X1 \DRAM_mem_reg[77][12]  ( .D(n6783), .CK(CLK), .QN(n35462) );
  DFF_X1 \DRAM_mem_reg[77][11]  ( .D(n6782), .CK(CLK), .QN(n35458) );
  DFF_X1 \DRAM_mem_reg[77][10]  ( .D(n6781), .CK(CLK), .QN(n35454) );
  DFF_X1 \DRAM_mem_reg[77][9]  ( .D(n6780), .CK(CLK), .QN(n35450) );
  DFF_X1 \DRAM_mem_reg[77][8]  ( .D(n6779), .CK(CLK), .QN(n35446) );
  DFF_X1 \DRAM_mem_reg[77][7]  ( .D(n6778), .CK(CLK), .QN(n35442) );
  DFF_X1 \DRAM_mem_reg[77][6]  ( .D(n6777), .CK(CLK), .QN(n35438) );
  DFF_X1 \DRAM_mem_reg[77][5]  ( .D(n6776), .CK(CLK), .QN(n35434) );
  DFF_X1 \DRAM_mem_reg[77][4]  ( .D(n6775), .CK(CLK), .QN(n35430) );
  DFF_X1 \DRAM_mem_reg[77][3]  ( .D(n6774), .CK(CLK), .QN(n35426) );
  DFF_X1 \DRAM_mem_reg[77][2]  ( .D(n6773), .CK(CLK), .QN(n35422) );
  DFF_X1 \DRAM_mem_reg[77][1]  ( .D(n6772), .CK(CLK), .QN(n35418) );
  DFF_X1 \DRAM_mem_reg[77][0]  ( .D(n6771), .CK(CLK), .QN(n35414) );
  DFF_X1 \DRAM_mem_reg[78][31]  ( .D(n6770), .CK(CLK), .Q(net253614), .QN(
        n37077) );
  DFF_X1 \DRAM_mem_reg[78][30]  ( .D(n6769), .CK(CLK), .Q(net253613), .QN(
        n37076) );
  DFF_X1 \DRAM_mem_reg[78][29]  ( .D(n6768), .CK(CLK), .Q(net253612), .QN(
        n37075) );
  DFF_X1 \DRAM_mem_reg[78][28]  ( .D(n6767), .CK(CLK), .Q(net253611), .QN(
        n37074) );
  DFF_X1 \DRAM_mem_reg[78][27]  ( .D(n6766), .CK(CLK), .Q(net253610), .QN(
        n37073) );
  DFF_X1 \DRAM_mem_reg[78][26]  ( .D(n6765), .CK(CLK), .Q(net253609), .QN(
        n37072) );
  DFF_X1 \DRAM_mem_reg[78][25]  ( .D(n6764), .CK(CLK), .Q(net253608), .QN(
        n37071) );
  DFF_X1 \DRAM_mem_reg[78][24]  ( .D(n6763), .CK(CLK), .Q(net253607), .QN(
        n37070) );
  DFF_X1 \DRAM_mem_reg[78][23]  ( .D(n6762), .CK(CLK), .Q(net253606), .QN(
        n37189) );
  DFF_X1 \DRAM_mem_reg[78][22]  ( .D(n6761), .CK(CLK), .Q(net253605), .QN(
        n37188) );
  DFF_X1 \DRAM_mem_reg[78][21]  ( .D(n6760), .CK(CLK), .Q(net253604), .QN(
        n37187) );
  DFF_X1 \DRAM_mem_reg[78][20]  ( .D(n6759), .CK(CLK), .Q(net253603), .QN(
        n37186) );
  DFF_X1 \DRAM_mem_reg[78][19]  ( .D(n6758), .CK(CLK), .Q(net253602), .QN(
        n37185) );
  DFF_X1 \DRAM_mem_reg[78][18]  ( .D(n6757), .CK(CLK), .Q(net253601), .QN(
        n37184) );
  DFF_X1 \DRAM_mem_reg[78][17]  ( .D(n6756), .CK(CLK), .Q(net253600), .QN(
        n37183) );
  DFF_X1 \DRAM_mem_reg[78][16]  ( .D(n6755), .CK(CLK), .Q(net253599), .QN(
        n37182) );
  DFF_X1 \DRAM_mem_reg[78][15]  ( .D(n6754), .CK(CLK), .Q(net253598), .QN(
        n37181) );
  DFF_X1 \DRAM_mem_reg[78][14]  ( .D(n6753), .CK(CLK), .Q(net253597), .QN(
        n37180) );
  DFF_X1 \DRAM_mem_reg[78][13]  ( .D(n6752), .CK(CLK), .Q(net253596), .QN(
        n37179) );
  DFF_X1 \DRAM_mem_reg[78][12]  ( .D(n6751), .CK(CLK), .Q(net253595), .QN(
        n37178) );
  DFF_X1 \DRAM_mem_reg[78][11]  ( .D(n6750), .CK(CLK), .Q(net253594), .QN(
        n37177) );
  DFF_X1 \DRAM_mem_reg[78][10]  ( .D(n6749), .CK(CLK), .Q(net253593), .QN(
        n37176) );
  DFF_X1 \DRAM_mem_reg[78][9]  ( .D(n6748), .CK(CLK), .Q(net253592), .QN(
        n37175) );
  DFF_X1 \DRAM_mem_reg[78][8]  ( .D(n6747), .CK(CLK), .Q(net253591), .QN(
        n37174) );
  DFF_X1 \DRAM_mem_reg[78][7]  ( .D(n6746), .CK(CLK), .Q(net253590), .QN(
        n37173) );
  DFF_X1 \DRAM_mem_reg[78][6]  ( .D(n6745), .CK(CLK), .Q(net253589), .QN(
        n37172) );
  DFF_X1 \DRAM_mem_reg[78][5]  ( .D(n6744), .CK(CLK), .Q(net253588), .QN(
        n37171) );
  DFF_X1 \DRAM_mem_reg[78][4]  ( .D(n6743), .CK(CLK), .Q(net253587), .QN(
        n37170) );
  DFF_X1 \DRAM_mem_reg[78][3]  ( .D(n6742), .CK(CLK), .Q(net253586), .QN(
        n37169) );
  DFF_X1 \DRAM_mem_reg[78][2]  ( .D(n6741), .CK(CLK), .Q(net253585), .QN(
        n37168) );
  DFF_X1 \DRAM_mem_reg[78][1]  ( .D(n6740), .CK(CLK), .Q(net253584), .QN(
        n37167) );
  DFF_X1 \DRAM_mem_reg[78][0]  ( .D(n6739), .CK(CLK), .Q(net253583), .QN(
        n37166) );
  DFF_X1 \DRAM_mem_reg[79][31]  ( .D(n6738), .CK(CLK), .Q(net253582), .QN(
        n37581) );
  DFF_X1 \Dout_reg[31]  ( .D(n6737), .CK(CLK), .Q(Dout[31]), .QN(n4145) );
  DFF_X1 \DRAM_mem_reg[79][30]  ( .D(n6736), .CK(CLK), .Q(net253581), .QN(
        n37580) );
  DFF_X1 \Dout_reg[30]  ( .D(n6735), .CK(CLK), .Q(Dout[30]), .QN(n4143) );
  DFF_X1 \DRAM_mem_reg[79][29]  ( .D(n6734), .CK(CLK), .Q(net253580), .QN(
        n37579) );
  DFF_X1 \Dout_reg[29]  ( .D(n6733), .CK(CLK), .Q(Dout[29]), .QN(n4141) );
  DFF_X1 \DRAM_mem_reg[79][28]  ( .D(n6732), .CK(CLK), .Q(net253579), .QN(
        n37578) );
  DFF_X1 \Dout_reg[28]  ( .D(n6731), .CK(CLK), .Q(Dout[28]), .QN(n4139) );
  DFF_X1 \DRAM_mem_reg[79][27]  ( .D(n6730), .CK(CLK), .Q(net253578), .QN(
        n37577) );
  DFF_X1 \Dout_reg[27]  ( .D(n6729), .CK(CLK), .Q(Dout[27]), .QN(n4137) );
  DFF_X1 \DRAM_mem_reg[79][26]  ( .D(n6728), .CK(CLK), .Q(net253577), .QN(
        n37576) );
  DFF_X1 \Dout_reg[26]  ( .D(n6727), .CK(CLK), .Q(Dout[26]), .QN(n4135) );
  DFF_X1 \DRAM_mem_reg[79][25]  ( .D(n6726), .CK(CLK), .Q(net253576), .QN(
        n37575) );
  DFF_X1 \Dout_reg[25]  ( .D(n6725), .CK(CLK), .Q(Dout[25]), .QN(n4133) );
  DFF_X1 \DRAM_mem_reg[79][24]  ( .D(n6724), .CK(CLK), .Q(net253575), .QN(
        n37574) );
  DFF_X1 \Dout_reg[24]  ( .D(n6723), .CK(CLK), .Q(Dout[24]), .QN(n4131) );
  DFF_X1 \DRAM_mem_reg[79][23]  ( .D(n6722), .CK(CLK), .Q(net253574), .QN(
        n37573) );
  DFF_X1 \Dout_reg[23]  ( .D(n6721), .CK(CLK), .Q(Dout[23]), .QN(n4129) );
  DFF_X1 \DRAM_mem_reg[79][22]  ( .D(n6720), .CK(CLK), .Q(net253573), .QN(
        n37572) );
  DFF_X1 \Dout_reg[22]  ( .D(n6719), .CK(CLK), .Q(Dout[22]), .QN(n4127) );
  DFF_X1 \DRAM_mem_reg[79][21]  ( .D(n6718), .CK(CLK), .Q(net253572), .QN(
        n37571) );
  DFF_X1 \Dout_reg[21]  ( .D(n6717), .CK(CLK), .Q(Dout[21]), .QN(n4125) );
  DFF_X1 \DRAM_mem_reg[79][20]  ( .D(n6716), .CK(CLK), .Q(net253571), .QN(
        n37570) );
  DFF_X1 \Dout_reg[20]  ( .D(n6715), .CK(CLK), .Q(Dout[20]), .QN(n4123) );
  DFF_X1 \DRAM_mem_reg[79][19]  ( .D(n6714), .CK(CLK), .Q(net253570), .QN(
        n37569) );
  DFF_X1 \Dout_reg[19]  ( .D(n6713), .CK(CLK), .Q(Dout[19]), .QN(n4121) );
  DFF_X1 \DRAM_mem_reg[79][18]  ( .D(n6712), .CK(CLK), .Q(net253569), .QN(
        n37568) );
  DFF_X1 \Dout_reg[18]  ( .D(n6711), .CK(CLK), .Q(Dout[18]), .QN(n4119) );
  DFF_X1 \DRAM_mem_reg[79][17]  ( .D(n6710), .CK(CLK), .Q(net253568), .QN(
        n37567) );
  DFF_X1 \Dout_reg[17]  ( .D(n6709), .CK(CLK), .Q(Dout[17]), .QN(n4117) );
  DFF_X1 \DRAM_mem_reg[79][16]  ( .D(n6708), .CK(CLK), .Q(net253567), .QN(
        n37566) );
  DFF_X1 \Dout_reg[16]  ( .D(n6707), .CK(CLK), .Q(Dout[16]), .QN(n4115) );
  DFF_X1 \DRAM_mem_reg[79][15]  ( .D(n6706), .CK(CLK), .Q(net253566), .QN(
        n37565) );
  DFF_X1 \Dout_reg[15]  ( .D(n6705), .CK(CLK), .Q(Dout[15]), .QN(n4113) );
  DFF_X1 \DRAM_mem_reg[79][14]  ( .D(n6704), .CK(CLK), .Q(net253565), .QN(
        n37564) );
  DFF_X1 \Dout_reg[14]  ( .D(n6703), .CK(CLK), .Q(Dout[14]), .QN(n4111) );
  DFF_X1 \DRAM_mem_reg[79][13]  ( .D(n6702), .CK(CLK), .Q(net253564), .QN(
        n37563) );
  DFF_X1 \Dout_reg[13]  ( .D(n6701), .CK(CLK), .Q(Dout[13]), .QN(n4109) );
  DFF_X1 \DRAM_mem_reg[79][12]  ( .D(n6700), .CK(CLK), .Q(net253563), .QN(
        n37562) );
  DFF_X1 \Dout_reg[12]  ( .D(n6699), .CK(CLK), .Q(Dout[12]), .QN(n4107) );
  DFF_X1 \DRAM_mem_reg[79][11]  ( .D(n6698), .CK(CLK), .Q(net253562), .QN(
        n37561) );
  DFF_X1 \Dout_reg[11]  ( .D(n6697), .CK(CLK), .Q(Dout[11]), .QN(n4105) );
  DFF_X1 \DRAM_mem_reg[79][10]  ( .D(n6696), .CK(CLK), .Q(net253561), .QN(
        n37560) );
  DFF_X1 \Dout_reg[10]  ( .D(n6695), .CK(CLK), .Q(Dout[10]), .QN(n4103) );
  DFF_X1 \DRAM_mem_reg[79][9]  ( .D(n6694), .CK(CLK), .Q(net253560), .QN(
        n37559) );
  DFF_X1 \Dout_reg[9]  ( .D(n6693), .CK(CLK), .Q(Dout[9]), .QN(n4101) );
  DFF_X1 \DRAM_mem_reg[79][8]  ( .D(n6692), .CK(CLK), .Q(net253559), .QN(
        n37558) );
  DFF_X1 \Dout_reg[8]  ( .D(n6691), .CK(CLK), .Q(Dout[8]), .QN(n4099) );
  DFF_X1 \DRAM_mem_reg[79][7]  ( .D(n6690), .CK(CLK), .Q(net253558), .QN(
        n37557) );
  DFF_X1 \Dout_reg[7]  ( .D(n6689), .CK(CLK), .Q(Dout[7]), .QN(n4097) );
  DFF_X1 \DRAM_mem_reg[79][6]  ( .D(n6688), .CK(CLK), .Q(net253557), .QN(
        n37556) );
  DFF_X1 \Dout_reg[6]  ( .D(n6687), .CK(CLK), .Q(Dout[6]), .QN(n4095) );
  DFF_X1 \DRAM_mem_reg[79][5]  ( .D(n6686), .CK(CLK), .Q(net253556), .QN(
        n37555) );
  DFF_X1 \Dout_reg[5]  ( .D(n6685), .CK(CLK), .Q(Dout[5]), .QN(n4093) );
  DFF_X1 \DRAM_mem_reg[79][4]  ( .D(n6684), .CK(CLK), .Q(net253555), .QN(
        n37554) );
  DFF_X1 \Dout_reg[4]  ( .D(n6683), .CK(CLK), .Q(Dout[4]), .QN(n4091) );
  DFF_X1 \DRAM_mem_reg[79][3]  ( .D(n6682), .CK(CLK), .Q(net253554), .QN(
        n37553) );
  DFF_X1 \Dout_reg[3]  ( .D(n6681), .CK(CLK), .Q(Dout[3]), .QN(n4089) );
  DFF_X1 \DRAM_mem_reg[79][2]  ( .D(n6680), .CK(CLK), .Q(net253553), .QN(
        n37552) );
  DFF_X1 \Dout_reg[2]  ( .D(n6679), .CK(CLK), .Q(Dout[2]), .QN(n4087) );
  DFF_X1 \DRAM_mem_reg[79][1]  ( .D(n6678), .CK(CLK), .Q(net253552), .QN(
        n37551) );
  DFF_X1 \Dout_reg[1]  ( .D(n6677), .CK(CLK), .Q(Dout[1]), .QN(n4085) );
  DFF_X1 \DRAM_mem_reg[79][0]  ( .D(n6676), .CK(CLK), .Q(net253551), .QN(
        n37550) );
  DFF_X1 \Dout_reg[0]  ( .D(n6675), .CK(CLK), .Q(Dout[0]), .QN(n4083) );
  NOR3_X2 U3 ( .A1(Addr[5]), .A2(Addr[6]), .A3(Addr[4]), .ZN(n9597) );
  NOR2_X2 U4 ( .A1(n9630), .A2(Addr[4]), .ZN(n9585) );
  NOR2_X2 U5 ( .A1(n9629), .A2(Addr[5]), .ZN(n9586) );
  OR3_X1 U6 ( .A1(n38911), .A2(WR_enable), .A3(n9631), .ZN(n35149) );
  INV_X1 U7 ( .A(n37977), .ZN(n37970) );
  INV_X1 U8 ( .A(n37989), .ZN(n37982) );
  INV_X1 U9 ( .A(n38010), .ZN(n38003) );
  INV_X1 U10 ( .A(n38031), .ZN(n38024) );
  INV_X1 U11 ( .A(n38043), .ZN(n38036) );
  INV_X1 U12 ( .A(n38052), .ZN(n38045) );
  INV_X1 U13 ( .A(n38064), .ZN(n38057) );
  INV_X1 U14 ( .A(n38085), .ZN(n38078) );
  INV_X1 U15 ( .A(n38097), .ZN(n38090) );
  INV_X1 U16 ( .A(n38118), .ZN(n38111) );
  INV_X1 U17 ( .A(n38139), .ZN(n38132) );
  INV_X1 U18 ( .A(n38151), .ZN(n38144) );
  INV_X1 U19 ( .A(n38172), .ZN(n38165) );
  INV_X1 U20 ( .A(n38184), .ZN(n38177) );
  INV_X1 U21 ( .A(n38205), .ZN(n38198) );
  INV_X1 U22 ( .A(n38226), .ZN(n38219) );
  INV_X1 U23 ( .A(n38238), .ZN(n38231) );
  INV_X1 U24 ( .A(n38259), .ZN(n38252) );
  INV_X1 U25 ( .A(n38280), .ZN(n38273) );
  INV_X1 U26 ( .A(n38292), .ZN(n38285) );
  INV_X1 U27 ( .A(n38313), .ZN(n38306) );
  INV_X1 U28 ( .A(n38325), .ZN(n38318) );
  INV_X1 U29 ( .A(n38346), .ZN(n38339) );
  INV_X1 U30 ( .A(n38367), .ZN(n38360) );
  INV_X1 U31 ( .A(n38379), .ZN(n38372) );
  INV_X1 U32 ( .A(n38400), .ZN(n38393) );
  INV_X1 U33 ( .A(n38421), .ZN(n38414) );
  INV_X1 U34 ( .A(n38433), .ZN(n38426) );
  INV_X1 U35 ( .A(n38454), .ZN(n38447) );
  INV_X1 U36 ( .A(n38475), .ZN(n38468) );
  INV_X1 U37 ( .A(n38493), .ZN(n38486) );
  INV_X1 U38 ( .A(n38505), .ZN(n38498) );
  INV_X1 U39 ( .A(n38553), .ZN(n38546) );
  INV_X1 U40 ( .A(n38565), .ZN(n38558) );
  INV_X1 U41 ( .A(n38613), .ZN(n38606) );
  INV_X1 U42 ( .A(n38625), .ZN(n38618) );
  INV_X1 U43 ( .A(n38673), .ZN(n38666) );
  INV_X1 U44 ( .A(n37998), .ZN(n37991) );
  INV_X1 U45 ( .A(n38019), .ZN(n38012) );
  INV_X1 U46 ( .A(n38073), .ZN(n38066) );
  INV_X1 U47 ( .A(n38106), .ZN(n38099) );
  INV_X1 U48 ( .A(n38127), .ZN(n38120) );
  INV_X1 U49 ( .A(n38160), .ZN(n38153) );
  INV_X1 U50 ( .A(n38193), .ZN(n38186) );
  INV_X1 U51 ( .A(n38214), .ZN(n38207) );
  INV_X1 U52 ( .A(n38247), .ZN(n38240) );
  INV_X1 U53 ( .A(n38268), .ZN(n38261) );
  INV_X1 U54 ( .A(n38301), .ZN(n38294) );
  INV_X1 U55 ( .A(n38334), .ZN(n38327) );
  INV_X1 U56 ( .A(n38355), .ZN(n38348) );
  INV_X1 U57 ( .A(n38388), .ZN(n38381) );
  INV_X1 U58 ( .A(n38409), .ZN(n38402) );
  INV_X1 U59 ( .A(n38442), .ZN(n38435) );
  INV_X1 U60 ( .A(n38463), .ZN(n38456) );
  INV_X1 U61 ( .A(n38909), .ZN(n38902) );
  BUF_X1 U62 ( .A(n37978), .Z(n37971) );
  BUF_X1 U63 ( .A(n37978), .Z(n37972) );
  BUF_X1 U64 ( .A(n37978), .Z(n37973) );
  BUF_X1 U65 ( .A(n37978), .Z(n37974) );
  BUF_X1 U66 ( .A(n37978), .Z(n37975) );
  BUF_X1 U67 ( .A(n37978), .Z(n37976) );
  BUF_X1 U68 ( .A(n37990), .Z(n37983) );
  BUF_X1 U69 ( .A(n37990), .Z(n37984) );
  BUF_X1 U70 ( .A(n37990), .Z(n37985) );
  BUF_X1 U71 ( .A(n37990), .Z(n37986) );
  BUF_X1 U72 ( .A(n37990), .Z(n37987) );
  BUF_X1 U73 ( .A(n37990), .Z(n37988) );
  BUF_X1 U74 ( .A(n38011), .Z(n38004) );
  BUF_X1 U75 ( .A(n38011), .Z(n38005) );
  BUF_X1 U76 ( .A(n38011), .Z(n38006) );
  BUF_X1 U77 ( .A(n38011), .Z(n38007) );
  BUF_X1 U78 ( .A(n38011), .Z(n38008) );
  BUF_X1 U79 ( .A(n38011), .Z(n38009) );
  BUF_X1 U80 ( .A(n38032), .Z(n38025) );
  BUF_X1 U81 ( .A(n38032), .Z(n38026) );
  BUF_X1 U82 ( .A(n38032), .Z(n38027) );
  BUF_X1 U83 ( .A(n38032), .Z(n38028) );
  BUF_X1 U84 ( .A(n38032), .Z(n38029) );
  BUF_X1 U85 ( .A(n38032), .Z(n38030) );
  BUF_X1 U86 ( .A(n38044), .Z(n38037) );
  BUF_X1 U87 ( .A(n38044), .Z(n38038) );
  BUF_X1 U88 ( .A(n38044), .Z(n38039) );
  BUF_X1 U89 ( .A(n38044), .Z(n38040) );
  BUF_X1 U90 ( .A(n38044), .Z(n38041) );
  BUF_X1 U91 ( .A(n38044), .Z(n38042) );
  BUF_X1 U92 ( .A(n38053), .Z(n38046) );
  BUF_X1 U93 ( .A(n38053), .Z(n38047) );
  BUF_X1 U94 ( .A(n38053), .Z(n38048) );
  BUF_X1 U95 ( .A(n38053), .Z(n38049) );
  BUF_X1 U96 ( .A(n38053), .Z(n38050) );
  BUF_X1 U97 ( .A(n38053), .Z(n38051) );
  BUF_X1 U98 ( .A(n38065), .Z(n38058) );
  BUF_X1 U99 ( .A(n38065), .Z(n38059) );
  BUF_X1 U100 ( .A(n38065), .Z(n38060) );
  BUF_X1 U101 ( .A(n38065), .Z(n38061) );
  BUF_X1 U102 ( .A(n38065), .Z(n38062) );
  BUF_X1 U103 ( .A(n38065), .Z(n38063) );
  BUF_X1 U104 ( .A(n38086), .Z(n38079) );
  BUF_X1 U105 ( .A(n38086), .Z(n38080) );
  BUF_X1 U106 ( .A(n38086), .Z(n38081) );
  BUF_X1 U107 ( .A(n38086), .Z(n38082) );
  BUF_X1 U108 ( .A(n38086), .Z(n38083) );
  BUF_X1 U109 ( .A(n38086), .Z(n38084) );
  BUF_X1 U110 ( .A(n38098), .Z(n38091) );
  BUF_X1 U111 ( .A(n38098), .Z(n38092) );
  BUF_X1 U112 ( .A(n38098), .Z(n38093) );
  BUF_X1 U113 ( .A(n38098), .Z(n38094) );
  BUF_X1 U114 ( .A(n38098), .Z(n38095) );
  BUF_X1 U115 ( .A(n38098), .Z(n38096) );
  BUF_X1 U116 ( .A(n38119), .Z(n38112) );
  BUF_X1 U117 ( .A(n38119), .Z(n38113) );
  BUF_X1 U118 ( .A(n38119), .Z(n38114) );
  BUF_X1 U119 ( .A(n38119), .Z(n38115) );
  BUF_X1 U120 ( .A(n38119), .Z(n38116) );
  BUF_X1 U121 ( .A(n38119), .Z(n38117) );
  BUF_X1 U122 ( .A(n38140), .Z(n38133) );
  BUF_X1 U123 ( .A(n38140), .Z(n38134) );
  BUF_X1 U124 ( .A(n38140), .Z(n38135) );
  BUF_X1 U125 ( .A(n38140), .Z(n38136) );
  BUF_X1 U126 ( .A(n38140), .Z(n38137) );
  BUF_X1 U127 ( .A(n38140), .Z(n38138) );
  BUF_X1 U128 ( .A(n38152), .Z(n38145) );
  BUF_X1 U129 ( .A(n38152), .Z(n38146) );
  BUF_X1 U130 ( .A(n38152), .Z(n38147) );
  BUF_X1 U131 ( .A(n38152), .Z(n38148) );
  BUF_X1 U132 ( .A(n38152), .Z(n38149) );
  BUF_X1 U133 ( .A(n38152), .Z(n38150) );
  BUF_X1 U134 ( .A(n38173), .Z(n38166) );
  BUF_X1 U135 ( .A(n38173), .Z(n38167) );
  BUF_X1 U136 ( .A(n38173), .Z(n38168) );
  BUF_X1 U137 ( .A(n38173), .Z(n38169) );
  BUF_X1 U138 ( .A(n38173), .Z(n38170) );
  BUF_X1 U139 ( .A(n38173), .Z(n38171) );
  BUF_X1 U140 ( .A(n38185), .Z(n38178) );
  BUF_X1 U141 ( .A(n38185), .Z(n38179) );
  BUF_X1 U142 ( .A(n38185), .Z(n38180) );
  BUF_X1 U143 ( .A(n38185), .Z(n38181) );
  BUF_X1 U144 ( .A(n38185), .Z(n38182) );
  BUF_X1 U145 ( .A(n38185), .Z(n38183) );
  BUF_X1 U146 ( .A(n38206), .Z(n38199) );
  BUF_X1 U147 ( .A(n38206), .Z(n38200) );
  BUF_X1 U148 ( .A(n38206), .Z(n38201) );
  BUF_X1 U149 ( .A(n38206), .Z(n38202) );
  BUF_X1 U150 ( .A(n38206), .Z(n38203) );
  BUF_X1 U151 ( .A(n38206), .Z(n38204) );
  BUF_X1 U152 ( .A(n38227), .Z(n38220) );
  BUF_X1 U153 ( .A(n38227), .Z(n38221) );
  BUF_X1 U154 ( .A(n38227), .Z(n38222) );
  BUF_X1 U155 ( .A(n38227), .Z(n38223) );
  BUF_X1 U156 ( .A(n38227), .Z(n38224) );
  BUF_X1 U157 ( .A(n38227), .Z(n38225) );
  BUF_X1 U158 ( .A(n38239), .Z(n38232) );
  BUF_X1 U159 ( .A(n38239), .Z(n38233) );
  BUF_X1 U160 ( .A(n38239), .Z(n38234) );
  BUF_X1 U161 ( .A(n38239), .Z(n38235) );
  BUF_X1 U162 ( .A(n38239), .Z(n38236) );
  BUF_X1 U163 ( .A(n38239), .Z(n38237) );
  BUF_X1 U164 ( .A(n38260), .Z(n38253) );
  BUF_X1 U165 ( .A(n38260), .Z(n38254) );
  BUF_X1 U166 ( .A(n38260), .Z(n38255) );
  BUF_X1 U167 ( .A(n38260), .Z(n38256) );
  BUF_X1 U168 ( .A(n38260), .Z(n38257) );
  BUF_X1 U169 ( .A(n38260), .Z(n38258) );
  BUF_X1 U170 ( .A(n38281), .Z(n38274) );
  BUF_X1 U171 ( .A(n38281), .Z(n38275) );
  BUF_X1 U172 ( .A(n38281), .Z(n38276) );
  BUF_X1 U173 ( .A(n38281), .Z(n38277) );
  BUF_X1 U174 ( .A(n38281), .Z(n38278) );
  BUF_X1 U175 ( .A(n38281), .Z(n38279) );
  BUF_X1 U176 ( .A(n38293), .Z(n38286) );
  BUF_X1 U177 ( .A(n38293), .Z(n38287) );
  BUF_X1 U178 ( .A(n38293), .Z(n38288) );
  BUF_X1 U179 ( .A(n38293), .Z(n38289) );
  BUF_X1 U180 ( .A(n38293), .Z(n38290) );
  BUF_X1 U181 ( .A(n38293), .Z(n38291) );
  BUF_X1 U182 ( .A(n38314), .Z(n38307) );
  BUF_X1 U183 ( .A(n38314), .Z(n38308) );
  BUF_X1 U184 ( .A(n38314), .Z(n38309) );
  BUF_X1 U185 ( .A(n38314), .Z(n38310) );
  BUF_X1 U186 ( .A(n38314), .Z(n38311) );
  BUF_X1 U187 ( .A(n38314), .Z(n38312) );
  BUF_X1 U188 ( .A(n38326), .Z(n38319) );
  BUF_X1 U189 ( .A(n38326), .Z(n38320) );
  BUF_X1 U190 ( .A(n38326), .Z(n38321) );
  BUF_X1 U191 ( .A(n38326), .Z(n38322) );
  BUF_X1 U192 ( .A(n38326), .Z(n38323) );
  BUF_X1 U193 ( .A(n38326), .Z(n38324) );
  BUF_X1 U194 ( .A(n38347), .Z(n38340) );
  BUF_X1 U195 ( .A(n38347), .Z(n38341) );
  BUF_X1 U196 ( .A(n38347), .Z(n38342) );
  BUF_X1 U197 ( .A(n38347), .Z(n38343) );
  BUF_X1 U198 ( .A(n38347), .Z(n38344) );
  BUF_X1 U199 ( .A(n38347), .Z(n38345) );
  BUF_X1 U200 ( .A(n38368), .Z(n38361) );
  BUF_X1 U201 ( .A(n38368), .Z(n38362) );
  BUF_X1 U202 ( .A(n38368), .Z(n38363) );
  BUF_X1 U203 ( .A(n38368), .Z(n38364) );
  BUF_X1 U204 ( .A(n38368), .Z(n38365) );
  BUF_X1 U205 ( .A(n38368), .Z(n38366) );
  BUF_X1 U206 ( .A(n38380), .Z(n38373) );
  BUF_X1 U207 ( .A(n38380), .Z(n38374) );
  BUF_X1 U208 ( .A(n38380), .Z(n38375) );
  BUF_X1 U209 ( .A(n38380), .Z(n38376) );
  BUF_X1 U210 ( .A(n38380), .Z(n38377) );
  BUF_X1 U211 ( .A(n38380), .Z(n38378) );
  BUF_X1 U212 ( .A(n38401), .Z(n38394) );
  BUF_X1 U213 ( .A(n38401), .Z(n38395) );
  BUF_X1 U214 ( .A(n38401), .Z(n38396) );
  BUF_X1 U215 ( .A(n38401), .Z(n38397) );
  BUF_X1 U216 ( .A(n38401), .Z(n38398) );
  BUF_X1 U217 ( .A(n38401), .Z(n38399) );
  BUF_X1 U218 ( .A(n38422), .Z(n38415) );
  BUF_X1 U219 ( .A(n38422), .Z(n38416) );
  BUF_X1 U220 ( .A(n38422), .Z(n38417) );
  BUF_X1 U221 ( .A(n38422), .Z(n38418) );
  BUF_X1 U222 ( .A(n38422), .Z(n38419) );
  BUF_X1 U223 ( .A(n38422), .Z(n38420) );
  BUF_X1 U224 ( .A(n38434), .Z(n38427) );
  BUF_X1 U225 ( .A(n38434), .Z(n38428) );
  BUF_X1 U226 ( .A(n38434), .Z(n38429) );
  BUF_X1 U227 ( .A(n38434), .Z(n38430) );
  BUF_X1 U228 ( .A(n38434), .Z(n38431) );
  BUF_X1 U229 ( .A(n38434), .Z(n38432) );
  BUF_X1 U230 ( .A(n38455), .Z(n38448) );
  BUF_X1 U231 ( .A(n38455), .Z(n38449) );
  BUF_X1 U232 ( .A(n38455), .Z(n38450) );
  BUF_X1 U233 ( .A(n38455), .Z(n38451) );
  BUF_X1 U234 ( .A(n38455), .Z(n38452) );
  BUF_X1 U235 ( .A(n38455), .Z(n38453) );
  BUF_X1 U236 ( .A(n38476), .Z(n38469) );
  BUF_X1 U237 ( .A(n38476), .Z(n38470) );
  BUF_X1 U238 ( .A(n38476), .Z(n38471) );
  BUF_X1 U239 ( .A(n38476), .Z(n38472) );
  BUF_X1 U240 ( .A(n38476), .Z(n38473) );
  BUF_X1 U241 ( .A(n38476), .Z(n38474) );
  BUF_X1 U242 ( .A(n38494), .Z(n38487) );
  BUF_X1 U243 ( .A(n38494), .Z(n38488) );
  BUF_X1 U244 ( .A(n38494), .Z(n38489) );
  BUF_X1 U245 ( .A(n38494), .Z(n38490) );
  BUF_X1 U246 ( .A(n38494), .Z(n38491) );
  BUF_X1 U247 ( .A(n38494), .Z(n38492) );
  BUF_X1 U248 ( .A(n37978), .Z(n37977) );
  BUF_X1 U249 ( .A(n37990), .Z(n37989) );
  BUF_X1 U250 ( .A(n38011), .Z(n38010) );
  BUF_X1 U251 ( .A(n38032), .Z(n38031) );
  BUF_X1 U252 ( .A(n38044), .Z(n38043) );
  BUF_X1 U253 ( .A(n38053), .Z(n38052) );
  BUF_X1 U254 ( .A(n38065), .Z(n38064) );
  BUF_X1 U255 ( .A(n38086), .Z(n38085) );
  BUF_X1 U256 ( .A(n38098), .Z(n38097) );
  BUF_X1 U257 ( .A(n38119), .Z(n38118) );
  BUF_X1 U258 ( .A(n38140), .Z(n38139) );
  BUF_X1 U259 ( .A(n38152), .Z(n38151) );
  BUF_X1 U260 ( .A(n38173), .Z(n38172) );
  BUF_X1 U261 ( .A(n38185), .Z(n38184) );
  BUF_X1 U262 ( .A(n38206), .Z(n38205) );
  BUF_X1 U263 ( .A(n38227), .Z(n38226) );
  BUF_X1 U264 ( .A(n38239), .Z(n38238) );
  BUF_X1 U265 ( .A(n38260), .Z(n38259) );
  BUF_X1 U266 ( .A(n38281), .Z(n38280) );
  BUF_X1 U267 ( .A(n38293), .Z(n38292) );
  BUF_X1 U268 ( .A(n38314), .Z(n38313) );
  BUF_X1 U269 ( .A(n38326), .Z(n38325) );
  BUF_X1 U270 ( .A(n38347), .Z(n38346) );
  BUF_X1 U271 ( .A(n38368), .Z(n38367) );
  BUF_X1 U272 ( .A(n38380), .Z(n38379) );
  BUF_X1 U273 ( .A(n38401), .Z(n38400) );
  BUF_X1 U274 ( .A(n38422), .Z(n38421) );
  BUF_X1 U275 ( .A(n38434), .Z(n38433) );
  BUF_X1 U276 ( .A(n38455), .Z(n38454) );
  BUF_X1 U277 ( .A(n38476), .Z(n38475) );
  BUF_X1 U278 ( .A(n38494), .Z(n38493) );
  BUF_X1 U279 ( .A(n5574), .Z(n37716) );
  BUF_X1 U280 ( .A(n5574), .Z(n37717) );
  BUF_X1 U281 ( .A(n5574), .Z(n37718) );
  INV_X1 U282 ( .A(n37804), .ZN(n37796) );
  INV_X1 U283 ( .A(n37804), .ZN(n37797) );
  INV_X1 U284 ( .A(n37812), .ZN(n37805) );
  INV_X1 U285 ( .A(n37824), .ZN(n37817) );
  INV_X1 U286 ( .A(n37836), .ZN(n37829) );
  INV_X1 U287 ( .A(n37848), .ZN(n37841) );
  INV_X1 U288 ( .A(n37857), .ZN(n37850) );
  INV_X1 U289 ( .A(n37866), .ZN(n37859) );
  INV_X1 U290 ( .A(n37878), .ZN(n37871) );
  INV_X1 U291 ( .A(n37890), .ZN(n37883) );
  INV_X1 U292 ( .A(n37902), .ZN(n37895) );
  INV_X1 U293 ( .A(n37911), .ZN(n37904) );
  INV_X1 U294 ( .A(n37920), .ZN(n37913) );
  INV_X1 U295 ( .A(n37932), .ZN(n37925) );
  INV_X1 U296 ( .A(n37944), .ZN(n37937) );
  INV_X1 U297 ( .A(n37956), .ZN(n37949) );
  INV_X1 U298 ( .A(n37965), .ZN(n37958) );
  INV_X1 U299 ( .A(n38517), .ZN(n38510) );
  INV_X1 U300 ( .A(n38529), .ZN(n38522) );
  INV_X1 U301 ( .A(n38541), .ZN(n38534) );
  INV_X1 U302 ( .A(n38577), .ZN(n38570) );
  INV_X1 U303 ( .A(n38589), .ZN(n38582) );
  INV_X1 U304 ( .A(n38601), .ZN(n38594) );
  INV_X1 U305 ( .A(n38637), .ZN(n38630) );
  INV_X1 U306 ( .A(n38649), .ZN(n38642) );
  INV_X1 U307 ( .A(n38661), .ZN(n38654) );
  INV_X1 U308 ( .A(n37795), .ZN(n37785) );
  INV_X1 U309 ( .A(n37795), .ZN(n37786) );
  BUF_X1 U310 ( .A(n37999), .Z(n37992) );
  BUF_X1 U311 ( .A(n37999), .Z(n37993) );
  BUF_X1 U312 ( .A(n37999), .Z(n37994) );
  BUF_X1 U313 ( .A(n37999), .Z(n37995) );
  BUF_X1 U314 ( .A(n37999), .Z(n37996) );
  BUF_X1 U315 ( .A(n37999), .Z(n37997) );
  BUF_X1 U316 ( .A(n38020), .Z(n38013) );
  BUF_X1 U317 ( .A(n38020), .Z(n38014) );
  BUF_X1 U318 ( .A(n38020), .Z(n38015) );
  BUF_X1 U319 ( .A(n38020), .Z(n38016) );
  BUF_X1 U320 ( .A(n38020), .Z(n38017) );
  BUF_X1 U321 ( .A(n38020), .Z(n38018) );
  BUF_X1 U322 ( .A(n38074), .Z(n38067) );
  BUF_X1 U323 ( .A(n38074), .Z(n38068) );
  BUF_X1 U324 ( .A(n38074), .Z(n38069) );
  BUF_X1 U325 ( .A(n38074), .Z(n38070) );
  BUF_X1 U326 ( .A(n38074), .Z(n38071) );
  BUF_X1 U327 ( .A(n38074), .Z(n38072) );
  BUF_X1 U328 ( .A(n38107), .Z(n38100) );
  BUF_X1 U329 ( .A(n38107), .Z(n38101) );
  BUF_X1 U330 ( .A(n38107), .Z(n38102) );
  BUF_X1 U331 ( .A(n38107), .Z(n38103) );
  BUF_X1 U332 ( .A(n38107), .Z(n38104) );
  BUF_X1 U333 ( .A(n38107), .Z(n38105) );
  BUF_X1 U334 ( .A(n38128), .Z(n38121) );
  BUF_X1 U335 ( .A(n38128), .Z(n38122) );
  BUF_X1 U336 ( .A(n38128), .Z(n38123) );
  BUF_X1 U337 ( .A(n38128), .Z(n38124) );
  BUF_X1 U338 ( .A(n38128), .Z(n38125) );
  BUF_X1 U339 ( .A(n38128), .Z(n38126) );
  BUF_X1 U340 ( .A(n38161), .Z(n38154) );
  BUF_X1 U341 ( .A(n38161), .Z(n38155) );
  BUF_X1 U342 ( .A(n38161), .Z(n38156) );
  BUF_X1 U343 ( .A(n38161), .Z(n38157) );
  BUF_X1 U344 ( .A(n38161), .Z(n38158) );
  BUF_X1 U345 ( .A(n38161), .Z(n38159) );
  BUF_X1 U346 ( .A(n38194), .Z(n38187) );
  BUF_X1 U347 ( .A(n38194), .Z(n38188) );
  BUF_X1 U348 ( .A(n38194), .Z(n38189) );
  BUF_X1 U349 ( .A(n38194), .Z(n38190) );
  BUF_X1 U350 ( .A(n38194), .Z(n38191) );
  BUF_X1 U351 ( .A(n38194), .Z(n38192) );
  BUF_X1 U352 ( .A(n38215), .Z(n38208) );
  BUF_X1 U353 ( .A(n38215), .Z(n38209) );
  BUF_X1 U354 ( .A(n38215), .Z(n38210) );
  BUF_X1 U355 ( .A(n38215), .Z(n38211) );
  BUF_X1 U356 ( .A(n38215), .Z(n38212) );
  BUF_X1 U357 ( .A(n38215), .Z(n38213) );
  BUF_X1 U358 ( .A(n38248), .Z(n38241) );
  BUF_X1 U359 ( .A(n38248), .Z(n38242) );
  BUF_X1 U360 ( .A(n38248), .Z(n38243) );
  BUF_X1 U361 ( .A(n38248), .Z(n38244) );
  BUF_X1 U362 ( .A(n38248), .Z(n38245) );
  BUF_X1 U363 ( .A(n38248), .Z(n38246) );
  BUF_X1 U364 ( .A(n38269), .Z(n38262) );
  BUF_X1 U365 ( .A(n38269), .Z(n38263) );
  BUF_X1 U366 ( .A(n38269), .Z(n38264) );
  BUF_X1 U367 ( .A(n38269), .Z(n38265) );
  BUF_X1 U368 ( .A(n38269), .Z(n38266) );
  BUF_X1 U369 ( .A(n38269), .Z(n38267) );
  BUF_X1 U370 ( .A(n38302), .Z(n38295) );
  BUF_X1 U371 ( .A(n38302), .Z(n38296) );
  BUF_X1 U372 ( .A(n38302), .Z(n38297) );
  BUF_X1 U373 ( .A(n38302), .Z(n38298) );
  BUF_X1 U374 ( .A(n38302), .Z(n38299) );
  BUF_X1 U375 ( .A(n38302), .Z(n38300) );
  BUF_X1 U376 ( .A(n38335), .Z(n38328) );
  BUF_X1 U377 ( .A(n38335), .Z(n38329) );
  BUF_X1 U378 ( .A(n38335), .Z(n38330) );
  BUF_X1 U379 ( .A(n38335), .Z(n38331) );
  BUF_X1 U380 ( .A(n38335), .Z(n38332) );
  BUF_X1 U381 ( .A(n38335), .Z(n38333) );
  BUF_X1 U382 ( .A(n38356), .Z(n38349) );
  BUF_X1 U383 ( .A(n38356), .Z(n38350) );
  BUF_X1 U384 ( .A(n38356), .Z(n38351) );
  BUF_X1 U385 ( .A(n38356), .Z(n38352) );
  BUF_X1 U386 ( .A(n38356), .Z(n38353) );
  BUF_X1 U387 ( .A(n38356), .Z(n38354) );
  BUF_X1 U388 ( .A(n38389), .Z(n38382) );
  BUF_X1 U389 ( .A(n38389), .Z(n38383) );
  BUF_X1 U390 ( .A(n38389), .Z(n38384) );
  BUF_X1 U391 ( .A(n38389), .Z(n38385) );
  BUF_X1 U392 ( .A(n38389), .Z(n38386) );
  BUF_X1 U393 ( .A(n38389), .Z(n38387) );
  BUF_X1 U394 ( .A(n38410), .Z(n38403) );
  BUF_X1 U395 ( .A(n38410), .Z(n38404) );
  BUF_X1 U396 ( .A(n38410), .Z(n38405) );
  BUF_X1 U397 ( .A(n38410), .Z(n38406) );
  BUF_X1 U398 ( .A(n38410), .Z(n38407) );
  BUF_X1 U399 ( .A(n38410), .Z(n38408) );
  BUF_X1 U400 ( .A(n38443), .Z(n38436) );
  BUF_X1 U401 ( .A(n38443), .Z(n38437) );
  BUF_X1 U402 ( .A(n38443), .Z(n38438) );
  BUF_X1 U403 ( .A(n38443), .Z(n38439) );
  BUF_X1 U404 ( .A(n38443), .Z(n38440) );
  BUF_X1 U405 ( .A(n38443), .Z(n38441) );
  BUF_X1 U406 ( .A(n38464), .Z(n38457) );
  BUF_X1 U407 ( .A(n38464), .Z(n38458) );
  BUF_X1 U408 ( .A(n38464), .Z(n38459) );
  BUF_X1 U409 ( .A(n38464), .Z(n38460) );
  BUF_X1 U410 ( .A(n38464), .Z(n38461) );
  BUF_X1 U411 ( .A(n38464), .Z(n38462) );
  BUF_X1 U412 ( .A(n38506), .Z(n38499) );
  BUF_X1 U413 ( .A(n38506), .Z(n38500) );
  BUF_X1 U414 ( .A(n38506), .Z(n38501) );
  BUF_X1 U415 ( .A(n38506), .Z(n38502) );
  BUF_X1 U416 ( .A(n38506), .Z(n38503) );
  BUF_X1 U417 ( .A(n38506), .Z(n38504) );
  BUF_X1 U418 ( .A(n38554), .Z(n38547) );
  BUF_X1 U419 ( .A(n38554), .Z(n38548) );
  BUF_X1 U420 ( .A(n38554), .Z(n38549) );
  BUF_X1 U421 ( .A(n38554), .Z(n38550) );
  BUF_X1 U422 ( .A(n38554), .Z(n38551) );
  BUF_X1 U423 ( .A(n38554), .Z(n38552) );
  BUF_X1 U424 ( .A(n38566), .Z(n38559) );
  BUF_X1 U425 ( .A(n38566), .Z(n38560) );
  BUF_X1 U426 ( .A(n38566), .Z(n38561) );
  BUF_X1 U427 ( .A(n38566), .Z(n38562) );
  BUF_X1 U428 ( .A(n38566), .Z(n38563) );
  BUF_X1 U429 ( .A(n38566), .Z(n38564) );
  BUF_X1 U430 ( .A(n38614), .Z(n38607) );
  BUF_X1 U431 ( .A(n38614), .Z(n38608) );
  BUF_X1 U432 ( .A(n38614), .Z(n38609) );
  BUF_X1 U433 ( .A(n38614), .Z(n38610) );
  BUF_X1 U434 ( .A(n38614), .Z(n38611) );
  BUF_X1 U435 ( .A(n38614), .Z(n38612) );
  BUF_X1 U436 ( .A(n38626), .Z(n38619) );
  BUF_X1 U437 ( .A(n38626), .Z(n38620) );
  BUF_X1 U438 ( .A(n38626), .Z(n38621) );
  BUF_X1 U439 ( .A(n38626), .Z(n38622) );
  BUF_X1 U440 ( .A(n38626), .Z(n38623) );
  BUF_X1 U441 ( .A(n38626), .Z(n38624) );
  BUF_X1 U442 ( .A(n38674), .Z(n38667) );
  BUF_X1 U443 ( .A(n38674), .Z(n38668) );
  BUF_X1 U444 ( .A(n38674), .Z(n38669) );
  BUF_X1 U445 ( .A(n38674), .Z(n38670) );
  BUF_X1 U446 ( .A(n38674), .Z(n38671) );
  BUF_X1 U447 ( .A(n38674), .Z(n38672) );
  BUF_X1 U448 ( .A(n38910), .Z(n38903) );
  BUF_X1 U449 ( .A(n38910), .Z(n38904) );
  BUF_X1 U450 ( .A(n38910), .Z(n38905) );
  BUF_X1 U451 ( .A(n38910), .Z(n38906) );
  BUF_X1 U452 ( .A(n38910), .Z(n38907) );
  BUF_X1 U453 ( .A(n38910), .Z(n38908) );
  BUF_X1 U454 ( .A(n37999), .Z(n37998) );
  BUF_X1 U455 ( .A(n38020), .Z(n38019) );
  BUF_X1 U456 ( .A(n38074), .Z(n38073) );
  BUF_X1 U457 ( .A(n38107), .Z(n38106) );
  BUF_X1 U458 ( .A(n38128), .Z(n38127) );
  BUF_X1 U459 ( .A(n38161), .Z(n38160) );
  BUF_X1 U460 ( .A(n38194), .Z(n38193) );
  BUF_X1 U461 ( .A(n38215), .Z(n38214) );
  BUF_X1 U462 ( .A(n38248), .Z(n38247) );
  BUF_X1 U463 ( .A(n38269), .Z(n38268) );
  BUF_X1 U464 ( .A(n38302), .Z(n38301) );
  BUF_X1 U465 ( .A(n38335), .Z(n38334) );
  BUF_X1 U466 ( .A(n38356), .Z(n38355) );
  BUF_X1 U467 ( .A(n38389), .Z(n38388) );
  BUF_X1 U468 ( .A(n38410), .Z(n38409) );
  BUF_X1 U469 ( .A(n38443), .Z(n38442) );
  BUF_X1 U470 ( .A(n38464), .Z(n38463) );
  BUF_X1 U471 ( .A(n38506), .Z(n38505) );
  BUF_X1 U472 ( .A(n38554), .Z(n38553) );
  BUF_X1 U473 ( .A(n38566), .Z(n38565) );
  BUF_X1 U474 ( .A(n38614), .Z(n38613) );
  BUF_X1 U475 ( .A(n38626), .Z(n38625) );
  BUF_X1 U476 ( .A(n38674), .Z(n38673) );
  BUF_X1 U477 ( .A(n38910), .Z(n38909) );
  INV_X1 U478 ( .A(n4843), .ZN(n38011) );
  OAI21_X1 U479 ( .B1(n38482), .B2(n38002), .A(n38920), .ZN(n4843) );
  INV_X1 U480 ( .A(n4668), .ZN(n38065) );
  OAI21_X1 U481 ( .B1(n38482), .B2(n38056), .A(n38920), .ZN(n4668) );
  INV_X1 U482 ( .A(n4493), .ZN(n38119) );
  OAI21_X1 U483 ( .B1(n38483), .B2(n38110), .A(n38920), .ZN(n4493) );
  INV_X1 U484 ( .A(n4388), .ZN(n38152) );
  OAI21_X1 U485 ( .B1(n38483), .B2(n38143), .A(n38919), .ZN(n4388) );
  INV_X1 U486 ( .A(n4213), .ZN(n38206) );
  OAI21_X1 U487 ( .B1(n38483), .B2(n38197), .A(n38919), .ZN(n4213) );
  INV_X1 U488 ( .A(n4006), .ZN(n38260) );
  OAI21_X1 U489 ( .B1(n38484), .B2(n38251), .A(n38919), .ZN(n4006) );
  INV_X1 U490 ( .A(n3831), .ZN(n38314) );
  OAI21_X1 U491 ( .B1(n38484), .B2(n38305), .A(n38918), .ZN(n3831) );
  INV_X1 U492 ( .A(n3726), .ZN(n38347) );
  OAI21_X1 U493 ( .B1(n38484), .B2(n38338), .A(n38918), .ZN(n3726) );
  INV_X1 U494 ( .A(n3551), .ZN(n38401) );
  OAI21_X1 U495 ( .B1(n38485), .B2(n38392), .A(n38918), .ZN(n3551) );
  INV_X1 U496 ( .A(n3376), .ZN(n38455) );
  OAI21_X1 U497 ( .B1(n38485), .B2(n38446), .A(n38917), .ZN(n3376) );
  INV_X1 U498 ( .A(n4703), .ZN(n38053) );
  OAI21_X1 U499 ( .B1(n38482), .B2(n4736), .A(n38920), .ZN(n4703) );
  INV_X1 U500 ( .A(n4948), .ZN(n37978) );
  OAI21_X1 U501 ( .B1(n38482), .B2(n37967), .A(n38917), .ZN(n4948) );
  INV_X1 U502 ( .A(n4913), .ZN(n37990) );
  OAI21_X1 U503 ( .B1(n38482), .B2(n37979), .A(n38919), .ZN(n4913) );
  INV_X1 U504 ( .A(n4773), .ZN(n38032) );
  OAI21_X1 U505 ( .B1(n38482), .B2(n38021), .A(n38920), .ZN(n4773) );
  INV_X1 U506 ( .A(n4738), .ZN(n38044) );
  OAI21_X1 U507 ( .B1(n38482), .B2(n38033), .A(n38920), .ZN(n4738) );
  INV_X1 U508 ( .A(n4598), .ZN(n38086) );
  OAI21_X1 U509 ( .B1(n38482), .B2(n38075), .A(n38920), .ZN(n4598) );
  INV_X1 U510 ( .A(n4563), .ZN(n38098) );
  OAI21_X1 U511 ( .B1(n38482), .B2(n38087), .A(n38920), .ZN(n4563) );
  INV_X1 U512 ( .A(n4423), .ZN(n38140) );
  OAI21_X1 U513 ( .B1(n38483), .B2(n38129), .A(n38919), .ZN(n4423) );
  INV_X1 U514 ( .A(n4318), .ZN(n38173) );
  OAI21_X1 U515 ( .B1(n38483), .B2(n38162), .A(n38919), .ZN(n4318) );
  INV_X1 U516 ( .A(n4283), .ZN(n38185) );
  OAI21_X1 U517 ( .B1(n38483), .B2(n38174), .A(n38919), .ZN(n4283) );
  INV_X1 U518 ( .A(n4140), .ZN(n38227) );
  OAI21_X1 U519 ( .B1(n38483), .B2(n38216), .A(n38919), .ZN(n4140) );
  INV_X1 U520 ( .A(n4076), .ZN(n38239) );
  OAI21_X1 U521 ( .B1(n38484), .B2(n38228), .A(n38919), .ZN(n4076) );
  INV_X1 U522 ( .A(n3936), .ZN(n38281) );
  OAI21_X1 U523 ( .B1(n38484), .B2(n38270), .A(n38918), .ZN(n3936) );
  INV_X1 U524 ( .A(n3901), .ZN(n38293) );
  OAI21_X1 U525 ( .B1(n38484), .B2(n38282), .A(n38918), .ZN(n3901) );
  INV_X1 U526 ( .A(n3796), .ZN(n38326) );
  OAI21_X1 U527 ( .B1(n38484), .B2(n38315), .A(n38918), .ZN(n3796) );
  INV_X1 U528 ( .A(n3656), .ZN(n38368) );
  OAI21_X1 U529 ( .B1(n38485), .B2(n38357), .A(n38918), .ZN(n3656) );
  INV_X1 U530 ( .A(n3621), .ZN(n38380) );
  OAI21_X1 U531 ( .B1(n38485), .B2(n38369), .A(n38918), .ZN(n3621) );
  INV_X1 U532 ( .A(n3481), .ZN(n38422) );
  OAI21_X1 U533 ( .B1(n38485), .B2(n38411), .A(n38917), .ZN(n3481) );
  INV_X1 U534 ( .A(n3446), .ZN(n38434) );
  OAI21_X1 U535 ( .B1(n38485), .B2(n38423), .A(n38917), .ZN(n3446) );
  INV_X1 U536 ( .A(n3306), .ZN(n38476) );
  OAI21_X1 U537 ( .B1(n38485), .B2(n38465), .A(n38917), .ZN(n3306) );
  INV_X1 U538 ( .A(n3270), .ZN(n38494) );
  OAI21_X1 U539 ( .B1(n38485), .B2(n38477), .A(n38917), .ZN(n3270) );
  BUF_X1 U540 ( .A(n5529), .Z(n37767) );
  BUF_X1 U541 ( .A(n5548), .Z(n37752) );
  BUF_X1 U542 ( .A(n5551), .Z(n37746) );
  BUF_X1 U543 ( .A(n5556), .Z(n37740) );
  BUF_X1 U544 ( .A(n5561), .Z(n37734) );
  BUF_X1 U545 ( .A(n5568), .Z(n37728) );
  BUF_X1 U546 ( .A(n5571), .Z(n37722) );
  BUF_X1 U547 ( .A(n5577), .Z(n37710) );
  BUF_X1 U548 ( .A(n5529), .Z(n37768) );
  BUF_X1 U549 ( .A(n5548), .Z(n37753) );
  BUF_X1 U550 ( .A(n5551), .Z(n37747) );
  BUF_X1 U551 ( .A(n5556), .Z(n37741) );
  BUF_X1 U552 ( .A(n5561), .Z(n37735) );
  BUF_X1 U553 ( .A(n5568), .Z(n37729) );
  BUF_X1 U554 ( .A(n5571), .Z(n37723) );
  BUF_X1 U555 ( .A(n5577), .Z(n37711) );
  BUF_X1 U556 ( .A(n4596), .Z(n38089) );
  BUF_X1 U557 ( .A(n4456), .Z(n38131) );
  BUF_X1 U558 ( .A(n4806), .Z(n38023) );
  BUF_X1 U559 ( .A(n4596), .Z(n38087) );
  BUF_X1 U560 ( .A(n4596), .Z(n38088) );
  BUF_X1 U561 ( .A(n4456), .Z(n38129) );
  BUF_X1 U562 ( .A(n4806), .Z(n38021) );
  BUF_X1 U563 ( .A(n4456), .Z(n38130) );
  BUF_X1 U564 ( .A(n4806), .Z(n38022) );
  BUF_X1 U565 ( .A(n5529), .Z(n37769) );
  BUF_X1 U566 ( .A(n5548), .Z(n37754) );
  BUF_X1 U567 ( .A(n5551), .Z(n37748) );
  BUF_X1 U568 ( .A(n5556), .Z(n37742) );
  BUF_X1 U569 ( .A(n5561), .Z(n37736) );
  BUF_X1 U570 ( .A(n5568), .Z(n37730) );
  BUF_X1 U571 ( .A(n5571), .Z(n37724) );
  BUF_X1 U572 ( .A(n5577), .Z(n37712) );
  BUF_X1 U573 ( .A(n5528), .Z(n37770) );
  BUF_X1 U574 ( .A(n5547), .Z(n37755) );
  BUF_X1 U575 ( .A(n5550), .Z(n37749) );
  BUF_X1 U576 ( .A(n5554), .Z(n37743) );
  BUF_X1 U577 ( .A(n5559), .Z(n37737) );
  BUF_X1 U578 ( .A(n5567), .Z(n37731) );
  BUF_X1 U579 ( .A(n5570), .Z(n37725) );
  BUF_X1 U580 ( .A(n5573), .Z(n37719) );
  BUF_X1 U581 ( .A(n5576), .Z(n37713) );
  BUF_X1 U582 ( .A(n5528), .Z(n37771) );
  BUF_X1 U583 ( .A(n5547), .Z(n37756) );
  BUF_X1 U584 ( .A(n5550), .Z(n37750) );
  BUF_X1 U585 ( .A(n5554), .Z(n37744) );
  BUF_X1 U586 ( .A(n5559), .Z(n37738) );
  BUF_X1 U587 ( .A(n5567), .Z(n37732) );
  BUF_X1 U588 ( .A(n5570), .Z(n37726) );
  BUF_X1 U589 ( .A(n5573), .Z(n37720) );
  BUF_X1 U590 ( .A(n5576), .Z(n37714) );
  BUF_X1 U591 ( .A(n5528), .Z(n37772) );
  BUF_X1 U592 ( .A(n5547), .Z(n37757) );
  BUF_X1 U593 ( .A(n5550), .Z(n37751) );
  BUF_X1 U594 ( .A(n5554), .Z(n37745) );
  BUF_X1 U595 ( .A(n5559), .Z(n37739) );
  BUF_X1 U596 ( .A(n5567), .Z(n37733) );
  BUF_X1 U597 ( .A(n5570), .Z(n37727) );
  BUF_X1 U598 ( .A(n5573), .Z(n37721) );
  BUF_X1 U599 ( .A(n5576), .Z(n37715) );
  INV_X1 U600 ( .A(n4736), .ZN(n5574) );
  INV_X1 U601 ( .A(n38913), .ZN(n38920) );
  INV_X1 U602 ( .A(n38913), .ZN(n38918) );
  INV_X1 U603 ( .A(n38913), .ZN(n38917) );
  INV_X1 U604 ( .A(n38913), .ZN(n38919) );
  INV_X1 U605 ( .A(n38913), .ZN(n38916) );
  BUF_X1 U606 ( .A(n38480), .Z(n38482) );
  BUF_X1 U607 ( .A(n38480), .Z(n38483) );
  BUF_X1 U608 ( .A(n38481), .Z(n38484) );
  BUF_X1 U609 ( .A(n38481), .Z(n38485) );
  BUF_X1 U610 ( .A(n5508), .Z(n37803) );
  BUF_X1 U611 ( .A(n5508), .Z(n37802) );
  BUF_X1 U612 ( .A(n5508), .Z(n37801) );
  BUF_X1 U613 ( .A(n5508), .Z(n37800) );
  BUF_X1 U614 ( .A(n5508), .Z(n37799) );
  BUF_X1 U615 ( .A(n5508), .Z(n37798) );
  BUF_X1 U616 ( .A(n38518), .Z(n38511) );
  BUF_X1 U617 ( .A(n38518), .Z(n38512) );
  BUF_X1 U618 ( .A(n38518), .Z(n38513) );
  BUF_X1 U619 ( .A(n38518), .Z(n38514) );
  BUF_X1 U620 ( .A(n38518), .Z(n38515) );
  BUF_X1 U621 ( .A(n38518), .Z(n38516) );
  BUF_X1 U622 ( .A(n38530), .Z(n38523) );
  BUF_X1 U623 ( .A(n38530), .Z(n38524) );
  BUF_X1 U624 ( .A(n38530), .Z(n38525) );
  BUF_X1 U625 ( .A(n38530), .Z(n38526) );
  BUF_X1 U626 ( .A(n38530), .Z(n38527) );
  BUF_X1 U627 ( .A(n38530), .Z(n38528) );
  BUF_X1 U628 ( .A(n38542), .Z(n38535) );
  BUF_X1 U629 ( .A(n38542), .Z(n38536) );
  BUF_X1 U630 ( .A(n38542), .Z(n38537) );
  BUF_X1 U631 ( .A(n38542), .Z(n38538) );
  BUF_X1 U632 ( .A(n38542), .Z(n38539) );
  BUF_X1 U633 ( .A(n38542), .Z(n38540) );
  BUF_X1 U634 ( .A(n38578), .Z(n38571) );
  BUF_X1 U635 ( .A(n38578), .Z(n38572) );
  BUF_X1 U636 ( .A(n38578), .Z(n38573) );
  BUF_X1 U637 ( .A(n38578), .Z(n38574) );
  BUF_X1 U638 ( .A(n38578), .Z(n38575) );
  BUF_X1 U639 ( .A(n38578), .Z(n38576) );
  BUF_X1 U640 ( .A(n38590), .Z(n38583) );
  BUF_X1 U641 ( .A(n38590), .Z(n38584) );
  BUF_X1 U642 ( .A(n38590), .Z(n38585) );
  BUF_X1 U643 ( .A(n38590), .Z(n38586) );
  BUF_X1 U644 ( .A(n38590), .Z(n38587) );
  BUF_X1 U645 ( .A(n38590), .Z(n38588) );
  BUF_X1 U646 ( .A(n38602), .Z(n38595) );
  BUF_X1 U647 ( .A(n38602), .Z(n38596) );
  BUF_X1 U648 ( .A(n38602), .Z(n38597) );
  BUF_X1 U649 ( .A(n38602), .Z(n38598) );
  BUF_X1 U650 ( .A(n38602), .Z(n38599) );
  BUF_X1 U651 ( .A(n38602), .Z(n38600) );
  BUF_X1 U652 ( .A(n38638), .Z(n38631) );
  BUF_X1 U653 ( .A(n38638), .Z(n38632) );
  BUF_X1 U654 ( .A(n38638), .Z(n38633) );
  BUF_X1 U655 ( .A(n38638), .Z(n38634) );
  BUF_X1 U656 ( .A(n38638), .Z(n38635) );
  BUF_X1 U657 ( .A(n38638), .Z(n38636) );
  BUF_X1 U658 ( .A(n38650), .Z(n38643) );
  BUF_X1 U659 ( .A(n38650), .Z(n38644) );
  BUF_X1 U660 ( .A(n38650), .Z(n38645) );
  BUF_X1 U661 ( .A(n38650), .Z(n38646) );
  BUF_X1 U662 ( .A(n38650), .Z(n38647) );
  BUF_X1 U663 ( .A(n38650), .Z(n38648) );
  BUF_X1 U664 ( .A(n38662), .Z(n38655) );
  BUF_X1 U665 ( .A(n38662), .Z(n38656) );
  BUF_X1 U666 ( .A(n38662), .Z(n38657) );
  BUF_X1 U667 ( .A(n38662), .Z(n38658) );
  BUF_X1 U668 ( .A(n38662), .Z(n38659) );
  BUF_X1 U669 ( .A(n38662), .Z(n38660) );
  BUF_X1 U670 ( .A(n37849), .Z(n37842) );
  BUF_X1 U671 ( .A(n37849), .Z(n37843) );
  BUF_X1 U672 ( .A(n37849), .Z(n37844) );
  BUF_X1 U673 ( .A(n37849), .Z(n37845) );
  BUF_X1 U674 ( .A(n37849), .Z(n37846) );
  BUF_X1 U675 ( .A(n37849), .Z(n37847) );
  BUF_X1 U676 ( .A(n37867), .Z(n37860) );
  BUF_X1 U677 ( .A(n37867), .Z(n37861) );
  BUF_X1 U678 ( .A(n37867), .Z(n37862) );
  BUF_X1 U679 ( .A(n37867), .Z(n37863) );
  BUF_X1 U680 ( .A(n37867), .Z(n37864) );
  BUF_X1 U681 ( .A(n37867), .Z(n37865) );
  BUF_X1 U682 ( .A(n37879), .Z(n37872) );
  BUF_X1 U683 ( .A(n37879), .Z(n37873) );
  BUF_X1 U684 ( .A(n37879), .Z(n37874) );
  BUF_X1 U685 ( .A(n37879), .Z(n37875) );
  BUF_X1 U686 ( .A(n37879), .Z(n37876) );
  BUF_X1 U687 ( .A(n37879), .Z(n37877) );
  BUF_X1 U688 ( .A(n37891), .Z(n37884) );
  BUF_X1 U689 ( .A(n37891), .Z(n37885) );
  BUF_X1 U690 ( .A(n37891), .Z(n37886) );
  BUF_X1 U691 ( .A(n37891), .Z(n37887) );
  BUF_X1 U692 ( .A(n37891), .Z(n37888) );
  BUF_X1 U693 ( .A(n37891), .Z(n37889) );
  BUF_X1 U694 ( .A(n37903), .Z(n37896) );
  BUF_X1 U695 ( .A(n37903), .Z(n37897) );
  BUF_X1 U696 ( .A(n37903), .Z(n37898) );
  BUF_X1 U697 ( .A(n37903), .Z(n37899) );
  BUF_X1 U698 ( .A(n37903), .Z(n37900) );
  BUF_X1 U699 ( .A(n37903), .Z(n37901) );
  BUF_X1 U700 ( .A(n37912), .Z(n37905) );
  BUF_X1 U701 ( .A(n37912), .Z(n37906) );
  BUF_X1 U702 ( .A(n37912), .Z(n37907) );
  BUF_X1 U703 ( .A(n37912), .Z(n37908) );
  BUF_X1 U704 ( .A(n37912), .Z(n37909) );
  BUF_X1 U705 ( .A(n37912), .Z(n37910) );
  BUF_X1 U706 ( .A(n37921), .Z(n37914) );
  BUF_X1 U707 ( .A(n37921), .Z(n37915) );
  BUF_X1 U708 ( .A(n37921), .Z(n37916) );
  BUF_X1 U709 ( .A(n37921), .Z(n37917) );
  BUF_X1 U710 ( .A(n37921), .Z(n37918) );
  BUF_X1 U711 ( .A(n37921), .Z(n37919) );
  BUF_X1 U712 ( .A(n37933), .Z(n37926) );
  BUF_X1 U713 ( .A(n37933), .Z(n37927) );
  BUF_X1 U714 ( .A(n37933), .Z(n37928) );
  BUF_X1 U715 ( .A(n37933), .Z(n37929) );
  BUF_X1 U716 ( .A(n37933), .Z(n37930) );
  BUF_X1 U717 ( .A(n37933), .Z(n37931) );
  BUF_X1 U718 ( .A(n37945), .Z(n37938) );
  BUF_X1 U719 ( .A(n37945), .Z(n37939) );
  BUF_X1 U720 ( .A(n37945), .Z(n37940) );
  BUF_X1 U721 ( .A(n37945), .Z(n37941) );
  BUF_X1 U722 ( .A(n37945), .Z(n37942) );
  BUF_X1 U723 ( .A(n37945), .Z(n37943) );
  BUF_X1 U724 ( .A(n37957), .Z(n37950) );
  BUF_X1 U725 ( .A(n37957), .Z(n37951) );
  BUF_X1 U726 ( .A(n37957), .Z(n37952) );
  BUF_X1 U727 ( .A(n37957), .Z(n37953) );
  BUF_X1 U728 ( .A(n37957), .Z(n37954) );
  BUF_X1 U729 ( .A(n37957), .Z(n37955) );
  BUF_X1 U730 ( .A(n37966), .Z(n37959) );
  BUF_X1 U731 ( .A(n37966), .Z(n37960) );
  BUF_X1 U732 ( .A(n37966), .Z(n37961) );
  BUF_X1 U733 ( .A(n37966), .Z(n37962) );
  BUF_X1 U734 ( .A(n37966), .Z(n37963) );
  BUF_X1 U735 ( .A(n37966), .Z(n37964) );
  BUF_X1 U736 ( .A(n37813), .Z(n37806) );
  BUF_X1 U737 ( .A(n37813), .Z(n37807) );
  BUF_X1 U738 ( .A(n37813), .Z(n37808) );
  BUF_X1 U739 ( .A(n37813), .Z(n37809) );
  BUF_X1 U740 ( .A(n37813), .Z(n37810) );
  BUF_X1 U741 ( .A(n37813), .Z(n37811) );
  BUF_X1 U742 ( .A(n37825), .Z(n37818) );
  BUF_X1 U743 ( .A(n37825), .Z(n37819) );
  BUF_X1 U744 ( .A(n37825), .Z(n37820) );
  BUF_X1 U745 ( .A(n37825), .Z(n37821) );
  BUF_X1 U746 ( .A(n37825), .Z(n37822) );
  BUF_X1 U747 ( .A(n37825), .Z(n37823) );
  BUF_X1 U748 ( .A(n37837), .Z(n37830) );
  BUF_X1 U749 ( .A(n37837), .Z(n37831) );
  BUF_X1 U750 ( .A(n37837), .Z(n37832) );
  BUF_X1 U751 ( .A(n37837), .Z(n37833) );
  BUF_X1 U752 ( .A(n37837), .Z(n37834) );
  BUF_X1 U753 ( .A(n37837), .Z(n37835) );
  BUF_X1 U754 ( .A(n37858), .Z(n37851) );
  BUF_X1 U755 ( .A(n37858), .Z(n37852) );
  BUF_X1 U756 ( .A(n37858), .Z(n37853) );
  BUF_X1 U757 ( .A(n37858), .Z(n37854) );
  BUF_X1 U758 ( .A(n37858), .Z(n37855) );
  BUF_X1 U759 ( .A(n37858), .Z(n37856) );
  BUF_X1 U760 ( .A(n5508), .Z(n37804) );
  BUF_X1 U761 ( .A(n38662), .Z(n38661) );
  BUF_X1 U762 ( .A(n38518), .Z(n38517) );
  BUF_X1 U763 ( .A(n38530), .Z(n38529) );
  BUF_X1 U764 ( .A(n38542), .Z(n38541) );
  BUF_X1 U765 ( .A(n38578), .Z(n38577) );
  BUF_X1 U766 ( .A(n38590), .Z(n38589) );
  BUF_X1 U767 ( .A(n38602), .Z(n38601) );
  BUF_X1 U768 ( .A(n38638), .Z(n38637) );
  BUF_X1 U769 ( .A(n38650), .Z(n38649) );
  BUF_X1 U770 ( .A(n37849), .Z(n37848) );
  BUF_X1 U771 ( .A(n37867), .Z(n37866) );
  BUF_X1 U772 ( .A(n37879), .Z(n37878) );
  BUF_X1 U773 ( .A(n37891), .Z(n37890) );
  BUF_X1 U774 ( .A(n37903), .Z(n37902) );
  BUF_X1 U775 ( .A(n37912), .Z(n37911) );
  BUF_X1 U776 ( .A(n37921), .Z(n37920) );
  BUF_X1 U777 ( .A(n37933), .Z(n37932) );
  BUF_X1 U778 ( .A(n37945), .Z(n37944) );
  BUF_X1 U779 ( .A(n37957), .Z(n37956) );
  BUF_X1 U780 ( .A(n37966), .Z(n37965) );
  BUF_X1 U781 ( .A(n37813), .Z(n37812) );
  BUF_X1 U782 ( .A(n37825), .Z(n37824) );
  BUF_X1 U783 ( .A(n37837), .Z(n37836) );
  BUF_X1 U784 ( .A(n37858), .Z(n37857) );
  BUF_X1 U785 ( .A(n35149), .Z(n37795) );
  BUF_X1 U786 ( .A(n37789), .Z(n37794) );
  BUF_X1 U787 ( .A(n37790), .Z(n37793) );
  BUF_X1 U788 ( .A(n35149), .Z(n37792) );
  BUF_X1 U789 ( .A(n35149), .Z(n37791) );
  BUF_X1 U790 ( .A(n35149), .Z(n37790) );
  BUF_X1 U791 ( .A(n35149), .Z(n37789) );
  BUF_X1 U792 ( .A(n35149), .Z(n37788) );
  BUF_X1 U793 ( .A(n35149), .Z(n37787) );
  INV_X1 U794 ( .A(n4878), .ZN(n37999) );
  OAI21_X1 U795 ( .B1(n38482), .B2(n4911), .A(n38920), .ZN(n4878) );
  INV_X1 U796 ( .A(n4808), .ZN(n38020) );
  OAI21_X1 U797 ( .B1(n38482), .B2(n4841), .A(n38920), .ZN(n4808) );
  INV_X1 U798 ( .A(n4633), .ZN(n38074) );
  OAI21_X1 U799 ( .B1(n38482), .B2(n4666), .A(n38920), .ZN(n4633) );
  INV_X1 U800 ( .A(n4528), .ZN(n38107) );
  OAI21_X1 U801 ( .B1(n38483), .B2(n4561), .A(n38920), .ZN(n4528) );
  INV_X1 U802 ( .A(n4458), .ZN(n38128) );
  OAI21_X1 U803 ( .B1(n38483), .B2(n4491), .A(n38920), .ZN(n4458) );
  INV_X1 U804 ( .A(n4353), .ZN(n38161) );
  OAI21_X1 U805 ( .B1(n38483), .B2(n4386), .A(n38919), .ZN(n4353) );
  INV_X1 U806 ( .A(n4248), .ZN(n38194) );
  OAI21_X1 U807 ( .B1(n38483), .B2(n4281), .A(n38919), .ZN(n4248) );
  INV_X1 U808 ( .A(n4178), .ZN(n38215) );
  OAI21_X1 U809 ( .B1(n38483), .B2(n4211), .A(n38919), .ZN(n4178) );
  INV_X1 U810 ( .A(n4041), .ZN(n38248) );
  OAI21_X1 U811 ( .B1(n38484), .B2(n4074), .A(n38919), .ZN(n4041) );
  INV_X1 U812 ( .A(n3971), .ZN(n38269) );
  OAI21_X1 U813 ( .B1(n38484), .B2(n4004), .A(n38918), .ZN(n3971) );
  INV_X1 U814 ( .A(n3866), .ZN(n38302) );
  OAI21_X1 U815 ( .B1(n38484), .B2(n3899), .A(n38918), .ZN(n3866) );
  INV_X1 U816 ( .A(n3761), .ZN(n38335) );
  OAI21_X1 U817 ( .B1(n38484), .B2(n3794), .A(n38918), .ZN(n3761) );
  INV_X1 U818 ( .A(n3691), .ZN(n38356) );
  OAI21_X1 U819 ( .B1(n38484), .B2(n3724), .A(n38918), .ZN(n3691) );
  INV_X1 U820 ( .A(n3586), .ZN(n38389) );
  OAI21_X1 U821 ( .B1(n38485), .B2(n3619), .A(n38918), .ZN(n3586) );
  INV_X1 U822 ( .A(n3516), .ZN(n38410) );
  OAI21_X1 U823 ( .B1(n38485), .B2(n3549), .A(n38917), .ZN(n3516) );
  INV_X1 U824 ( .A(n3411), .ZN(n38443) );
  OAI21_X1 U825 ( .B1(n38485), .B2(n3444), .A(n38917), .ZN(n3411) );
  INV_X1 U826 ( .A(n3341), .ZN(n38464) );
  OAI21_X1 U827 ( .B1(n38485), .B2(n3374), .A(n38917), .ZN(n3341) );
  INV_X1 U828 ( .A(n3236), .ZN(n38506) );
  OAI21_X1 U829 ( .B1(n38912), .B2(n38495), .A(n2741), .ZN(n3236) );
  INV_X1 U830 ( .A(n3096), .ZN(n38554) );
  OAI21_X1 U831 ( .B1(n38912), .B2(n38543), .A(n2741), .ZN(n3096) );
  INV_X1 U832 ( .A(n3061), .ZN(n38566) );
  OAI21_X1 U833 ( .B1(n38912), .B2(n38555), .A(n2741), .ZN(n3061) );
  INV_X1 U834 ( .A(n2921), .ZN(n38614) );
  OAI21_X1 U835 ( .B1(n38912), .B2(n38603), .A(n2741), .ZN(n2921) );
  INV_X1 U836 ( .A(n2886), .ZN(n38626) );
  OAI21_X1 U837 ( .B1(n38911), .B2(n38615), .A(n2741), .ZN(n2886) );
  INV_X1 U838 ( .A(n2744), .ZN(n38674) );
  OAI21_X1 U839 ( .B1(n38911), .B2(n38663), .A(n2741), .ZN(n2744) );
  INV_X1 U840 ( .A(n2676), .ZN(n38910) );
  OAI21_X1 U841 ( .B1(n38911), .B2(n38675), .A(n2741), .ZN(n2676) );
  BUF_X1 U842 ( .A(n5523), .Z(n37779) );
  BUF_X1 U843 ( .A(n5526), .Z(n37773) );
  BUF_X1 U844 ( .A(n5532), .Z(n37761) );
  BUF_X1 U845 ( .A(n5540), .Z(n37758) );
  BUF_X1 U846 ( .A(n5523), .Z(n37780) );
  BUF_X1 U847 ( .A(n5526), .Z(n37774) );
  BUF_X1 U848 ( .A(n5532), .Z(n37762) );
  BUF_X1 U849 ( .A(n5540), .Z(n37759) );
  BUF_X1 U850 ( .A(n3128), .Z(n38543) );
  BUF_X1 U851 ( .A(n2953), .Z(n38603) );
  BUF_X1 U852 ( .A(n2776), .Z(n38663) );
  BUF_X1 U853 ( .A(n2953), .Z(n38604) );
  BUF_X1 U854 ( .A(n2776), .Z(n38664) );
  BUF_X1 U855 ( .A(n3128), .Z(n38544) );
  BUF_X1 U856 ( .A(n4526), .Z(n38110) );
  BUF_X1 U857 ( .A(n3864), .Z(n38305) );
  BUF_X1 U858 ( .A(n3023), .Z(n38581) );
  BUF_X1 U859 ( .A(n2848), .Z(n38641) );
  BUF_X1 U860 ( .A(n3198), .Z(n38521) );
  BUF_X1 U861 ( .A(n4876), .Z(n38002) );
  BUF_X1 U862 ( .A(n4246), .Z(n38197) );
  BUF_X1 U863 ( .A(n4421), .Z(n38143) );
  BUF_X1 U864 ( .A(n3759), .Z(n38338) );
  BUF_X1 U865 ( .A(n4039), .Z(n38251) );
  BUF_X1 U866 ( .A(n3409), .Z(n38446) );
  BUF_X1 U867 ( .A(n3584), .Z(n38392) );
  BUF_X1 U868 ( .A(n4701), .Z(n38056) );
  BUF_X1 U869 ( .A(n3934), .Z(n38284) );
  BUF_X1 U870 ( .A(n3304), .Z(n38479) );
  BUF_X1 U871 ( .A(n3058), .Z(n38569) );
  BUF_X1 U872 ( .A(n2883), .Z(n38629) );
  BUF_X1 U873 ( .A(n3233), .Z(n38509) );
  BUF_X1 U874 ( .A(n4316), .Z(n38176) );
  BUF_X1 U875 ( .A(n3654), .Z(n38371) );
  BUF_X1 U876 ( .A(n3829), .Z(n38317) );
  BUF_X1 U877 ( .A(n4946), .Z(n37981) );
  BUF_X1 U878 ( .A(n3479), .Z(n38425) );
  BUF_X1 U879 ( .A(n4771), .Z(n38035) );
  BUF_X1 U880 ( .A(n4136), .Z(n38230) );
  BUF_X1 U881 ( .A(n4526), .Z(n38108) );
  BUF_X1 U882 ( .A(n3864), .Z(n38303) );
  BUF_X1 U883 ( .A(n3023), .Z(n38579) );
  BUF_X1 U884 ( .A(n2848), .Z(n38639) );
  BUF_X1 U885 ( .A(n3198), .Z(n38519) );
  BUF_X1 U886 ( .A(n4876), .Z(n38000) );
  BUF_X1 U887 ( .A(n4246), .Z(n38195) );
  BUF_X1 U888 ( .A(n4421), .Z(n38141) );
  BUF_X1 U889 ( .A(n3759), .Z(n38336) );
  BUF_X1 U890 ( .A(n4039), .Z(n38249) );
  BUF_X1 U891 ( .A(n3409), .Z(n38444) );
  BUF_X1 U892 ( .A(n3584), .Z(n38390) );
  BUF_X1 U893 ( .A(n4701), .Z(n38054) );
  BUF_X1 U894 ( .A(n4526), .Z(n38109) );
  BUF_X1 U895 ( .A(n3864), .Z(n38304) );
  BUF_X1 U896 ( .A(n3023), .Z(n38580) );
  BUF_X1 U897 ( .A(n2848), .Z(n38640) );
  BUF_X1 U898 ( .A(n3198), .Z(n38520) );
  BUF_X1 U899 ( .A(n4876), .Z(n38001) );
  BUF_X1 U900 ( .A(n4246), .Z(n38196) );
  BUF_X1 U901 ( .A(n4421), .Z(n38142) );
  BUF_X1 U902 ( .A(n3759), .Z(n38337) );
  BUF_X1 U903 ( .A(n4039), .Z(n38250) );
  BUF_X1 U904 ( .A(n3409), .Z(n38445) );
  BUF_X1 U905 ( .A(n3584), .Z(n38391) );
  BUF_X1 U906 ( .A(n4701), .Z(n38055) );
  BUF_X1 U907 ( .A(n3339), .Z(n38467) );
  BUF_X1 U908 ( .A(n2988), .Z(n38593) );
  BUF_X1 U909 ( .A(n3163), .Z(n38533) );
  BUF_X1 U910 ( .A(n3689), .Z(n38359) );
  BUF_X1 U911 ( .A(n4981), .Z(n37969) );
  BUF_X1 U912 ( .A(n4351), .Z(n38164) );
  BUF_X1 U913 ( .A(n4631), .Z(n38077) );
  BUF_X1 U914 ( .A(n3969), .Z(n38272) );
  BUF_X1 U915 ( .A(n4176), .Z(n38218) );
  BUF_X1 U916 ( .A(n3514), .Z(n38413) );
  BUF_X1 U917 ( .A(n2918), .Z(n38617) );
  BUF_X1 U918 ( .A(n2740), .Z(n38677) );
  BUF_X1 U919 ( .A(n3268), .Z(n38497) );
  BUF_X1 U920 ( .A(n3093), .Z(n38557) );
  BUF_X1 U921 ( .A(n3934), .Z(n38282) );
  BUF_X1 U922 ( .A(n3304), .Z(n38477) );
  BUF_X1 U923 ( .A(n3058), .Z(n38567) );
  BUF_X1 U924 ( .A(n2883), .Z(n38627) );
  BUF_X1 U925 ( .A(n3233), .Z(n38507) );
  BUF_X1 U926 ( .A(n4316), .Z(n38174) );
  BUF_X1 U927 ( .A(n3654), .Z(n38369) );
  BUF_X1 U928 ( .A(n3829), .Z(n38315) );
  BUF_X1 U929 ( .A(n4946), .Z(n37979) );
  BUF_X1 U930 ( .A(n3479), .Z(n38423) );
  BUF_X1 U931 ( .A(n4771), .Z(n38033) );
  BUF_X1 U932 ( .A(n4136), .Z(n38228) );
  BUF_X1 U933 ( .A(n3934), .Z(n38283) );
  BUF_X1 U934 ( .A(n3304), .Z(n38478) );
  BUF_X1 U935 ( .A(n3058), .Z(n38568) );
  BUF_X1 U936 ( .A(n2883), .Z(n38628) );
  BUF_X1 U937 ( .A(n3233), .Z(n38508) );
  BUF_X1 U938 ( .A(n4316), .Z(n38175) );
  BUF_X1 U939 ( .A(n3654), .Z(n38370) );
  BUF_X1 U940 ( .A(n3829), .Z(n38316) );
  BUF_X1 U941 ( .A(n4946), .Z(n37980) );
  BUF_X1 U942 ( .A(n3479), .Z(n38424) );
  BUF_X1 U943 ( .A(n4771), .Z(n38034) );
  BUF_X1 U944 ( .A(n4136), .Z(n38229) );
  BUF_X1 U945 ( .A(n2811), .Z(n38653) );
  BUF_X1 U946 ( .A(n3339), .Z(n38465) );
  BUF_X1 U947 ( .A(n2988), .Z(n38591) );
  BUF_X1 U948 ( .A(n3163), .Z(n38531) );
  BUF_X1 U949 ( .A(n3689), .Z(n38357) );
  BUF_X1 U950 ( .A(n4981), .Z(n37967) );
  BUF_X1 U951 ( .A(n4351), .Z(n38162) );
  BUF_X1 U952 ( .A(n4631), .Z(n38075) );
  BUF_X1 U953 ( .A(n3969), .Z(n38270) );
  BUF_X1 U954 ( .A(n4176), .Z(n38216) );
  BUF_X1 U955 ( .A(n3514), .Z(n38411) );
  BUF_X1 U956 ( .A(n3268), .Z(n38495) );
  BUF_X1 U957 ( .A(n3093), .Z(n38555) );
  BUF_X1 U958 ( .A(n2918), .Z(n38615) );
  BUF_X1 U959 ( .A(n2740), .Z(n38675) );
  BUF_X1 U960 ( .A(n2811), .Z(n38651) );
  BUF_X1 U961 ( .A(n3339), .Z(n38466) );
  BUF_X1 U962 ( .A(n2988), .Z(n38592) );
  BUF_X1 U963 ( .A(n3163), .Z(n38532) );
  BUF_X1 U964 ( .A(n3689), .Z(n38358) );
  BUF_X1 U965 ( .A(n4981), .Z(n37968) );
  BUF_X1 U966 ( .A(n4351), .Z(n38163) );
  BUF_X1 U967 ( .A(n4631), .Z(n38076) );
  BUF_X1 U968 ( .A(n3969), .Z(n38271) );
  BUF_X1 U969 ( .A(n4176), .Z(n38217) );
  BUF_X1 U970 ( .A(n3514), .Z(n38412) );
  BUF_X1 U971 ( .A(n2811), .Z(n38652) );
  BUF_X1 U972 ( .A(n2918), .Z(n38616) );
  BUF_X1 U973 ( .A(n2740), .Z(n38676) );
  BUF_X1 U974 ( .A(n3268), .Z(n38496) );
  BUF_X1 U975 ( .A(n3093), .Z(n38556) );
  BUF_X1 U976 ( .A(n5523), .Z(n37781) );
  BUF_X1 U977 ( .A(n5526), .Z(n37775) );
  BUF_X1 U978 ( .A(n5532), .Z(n37763) );
  BUF_X1 U979 ( .A(n5540), .Z(n37760) );
  BUF_X1 U980 ( .A(n5522), .Z(n37782) );
  BUF_X1 U981 ( .A(n5525), .Z(n37776) );
  BUF_X1 U982 ( .A(n5531), .Z(n37764) );
  BUF_X1 U983 ( .A(n5522), .Z(n37783) );
  BUF_X1 U984 ( .A(n5525), .Z(n37777) );
  BUF_X1 U985 ( .A(n5531), .Z(n37765) );
  BUF_X1 U986 ( .A(n5522), .Z(n37784) );
  BUF_X1 U987 ( .A(n5525), .Z(n37778) );
  BUF_X1 U988 ( .A(n5531), .Z(n37766) );
  NAND2_X1 U989 ( .A1(n9583), .A2(n9589), .ZN(n4456) );
  NAND2_X1 U990 ( .A1(n9583), .A2(n9574), .ZN(n4806) );
  NAND2_X1 U991 ( .A1(n9583), .A2(n9581), .ZN(n4596) );
  NAND2_X1 U992 ( .A1(n9583), .A2(n9578), .ZN(n4736) );
  BUF_X1 U993 ( .A(n2953), .Z(n38605) );
  BUF_X1 U994 ( .A(n2776), .Z(n38665) );
  BUF_X1 U995 ( .A(n3128), .Z(n38545) );
  INV_X1 U996 ( .A(n3899), .ZN(n5529) );
  INV_X1 U997 ( .A(n4491), .ZN(n5528) );
  INV_X1 U998 ( .A(n4281), .ZN(n5548) );
  INV_X1 U999 ( .A(n4841), .ZN(n5547) );
  INV_X1 U1000 ( .A(n3619), .ZN(n5551) );
  INV_X1 U1001 ( .A(n4211), .ZN(n5550) );
  INV_X1 U1002 ( .A(n3794), .ZN(n5556) );
  INV_X1 U1003 ( .A(n4386), .ZN(n5554) );
  INV_X1 U1004 ( .A(n4911), .ZN(n5561) );
  INV_X1 U1005 ( .A(n3724), .ZN(n5559) );
  INV_X1 U1006 ( .A(n3444), .ZN(n5568) );
  INV_X1 U1007 ( .A(n4004), .ZN(n5567) );
  INV_X1 U1008 ( .A(n4561), .ZN(n5571) );
  INV_X1 U1009 ( .A(n3374), .ZN(n5570) );
  INV_X1 U1010 ( .A(n3549), .ZN(n5573) );
  INV_X1 U1011 ( .A(n4074), .ZN(n5577) );
  INV_X1 U1012 ( .A(n4666), .ZN(n5576) );
  OAI222_X1 U1013 ( .A1(n37892), .A2(n35662), .B1(n37868), .B2(n35150), .C1(
        n37882), .C2(n36174), .ZN(n5842) );
  OAI222_X1 U1014 ( .A1(n38465), .A2(n35686), .B1(n38282), .B2(n35166), .C1(
        n38110), .C2(n36190), .ZN(n5843) );
  OAI222_X1 U1015 ( .A1(n38129), .A2(n35678), .B1(n38477), .B2(n35174), .C1(
        n38305), .C2(n36198), .ZN(n5844) );
  OAI222_X1 U1016 ( .A1(n38653), .A2(n35702), .B1(n38627), .B2(n35190), .C1(
        n38641), .C2(n36214), .ZN(n5850) );
  OAI222_X1 U1017 ( .A1(n37946), .A2(n35670), .B1(n37922), .B2(n35158), .C1(
        n37936), .C2(n36182), .ZN(n5851) );
  OAI222_X1 U1018 ( .A1(n38531), .A2(n35694), .B1(n38507), .B2(n35182), .C1(
        n38521), .C2(n36206), .ZN(n5852) );
  OAI222_X1 U1019 ( .A1(n37892), .A2(n35663), .B1(n37868), .B2(n35151), .C1(
        n37882), .C2(n36175), .ZN(n5800) );
  OAI222_X1 U1020 ( .A1(n38465), .A2(n35687), .B1(n38282), .B2(n35167), .C1(
        n38110), .C2(n36191), .ZN(n5801) );
  OAI222_X1 U1021 ( .A1(n38129), .A2(n35679), .B1(n38477), .B2(n35175), .C1(
        n38305), .C2(n36199), .ZN(n5802) );
  OAI222_X1 U1022 ( .A1(n38653), .A2(n35703), .B1(n38627), .B2(n35191), .C1(
        n38641), .C2(n36215), .ZN(n5808) );
  OAI222_X1 U1023 ( .A1(n37946), .A2(n35671), .B1(n37922), .B2(n35159), .C1(
        n37936), .C2(n36183), .ZN(n5809) );
  OAI222_X1 U1024 ( .A1(n38531), .A2(n35695), .B1(n38507), .B2(n35183), .C1(
        n38521), .C2(n36207), .ZN(n5810) );
  OAI222_X1 U1025 ( .A1(n37892), .A2(n35664), .B1(n37868), .B2(n35152), .C1(
        n37882), .C2(n36176), .ZN(n5758) );
  OAI222_X1 U1026 ( .A1(n38465), .A2(n35688), .B1(n38282), .B2(n35168), .C1(
        n38110), .C2(n36192), .ZN(n5759) );
  OAI222_X1 U1027 ( .A1(n38129), .A2(n35680), .B1(n38477), .B2(n35176), .C1(
        n38305), .C2(n36200), .ZN(n5760) );
  OAI222_X1 U1028 ( .A1(n38653), .A2(n35704), .B1(n38627), .B2(n35192), .C1(
        n38641), .C2(n36216), .ZN(n5766) );
  OAI222_X1 U1029 ( .A1(n37946), .A2(n35672), .B1(n37922), .B2(n35160), .C1(
        n37936), .C2(n36184), .ZN(n5767) );
  OAI222_X1 U1030 ( .A1(n38531), .A2(n35696), .B1(n38507), .B2(n35184), .C1(
        n38521), .C2(n36208), .ZN(n5768) );
  OAI222_X1 U1031 ( .A1(n37892), .A2(n35665), .B1(n37868), .B2(n35153), .C1(
        n37882), .C2(n36177), .ZN(n5716) );
  OAI222_X1 U1032 ( .A1(n38465), .A2(n35689), .B1(n38282), .B2(n35169), .C1(
        n38110), .C2(n36193), .ZN(n5717) );
  OAI222_X1 U1033 ( .A1(n38129), .A2(n35681), .B1(n38477), .B2(n35177), .C1(
        n38305), .C2(n36201), .ZN(n5718) );
  OAI222_X1 U1034 ( .A1(n38653), .A2(n35705), .B1(n38627), .B2(n35193), .C1(
        n38641), .C2(n36217), .ZN(n5724) );
  OAI222_X1 U1035 ( .A1(n37946), .A2(n35673), .B1(n37922), .B2(n35161), .C1(
        n37936), .C2(n36185), .ZN(n5725) );
  OAI222_X1 U1036 ( .A1(n38531), .A2(n35697), .B1(n38507), .B2(n35185), .C1(
        n38521), .C2(n36209), .ZN(n5726) );
  OAI222_X1 U1037 ( .A1(n37892), .A2(n35666), .B1(n37868), .B2(n35154), .C1(
        n37882), .C2(n36178), .ZN(n5674) );
  OAI222_X1 U1038 ( .A1(n38465), .A2(n35690), .B1(n38282), .B2(n35170), .C1(
        n38110), .C2(n36194), .ZN(n5675) );
  OAI222_X1 U1039 ( .A1(n38129), .A2(n35682), .B1(n38477), .B2(n35178), .C1(
        n38305), .C2(n36202), .ZN(n5676) );
  OAI222_X1 U1040 ( .A1(n38653), .A2(n35706), .B1(n38627), .B2(n35194), .C1(
        n38641), .C2(n36218), .ZN(n5682) );
  OAI222_X1 U1041 ( .A1(n37946), .A2(n35674), .B1(n37922), .B2(n35162), .C1(
        n37936), .C2(n36186), .ZN(n5683) );
  OAI222_X1 U1042 ( .A1(n38531), .A2(n35698), .B1(n38507), .B2(n35186), .C1(
        n38521), .C2(n36210), .ZN(n5684) );
  OAI222_X1 U1043 ( .A1(n37892), .A2(n35667), .B1(n37868), .B2(n35155), .C1(
        n37882), .C2(n36179), .ZN(n5632) );
  OAI222_X1 U1044 ( .A1(n38465), .A2(n35691), .B1(n38282), .B2(n35171), .C1(
        n38110), .C2(n36195), .ZN(n5633) );
  OAI222_X1 U1045 ( .A1(n38129), .A2(n35683), .B1(n38477), .B2(n35179), .C1(
        n38305), .C2(n36203), .ZN(n5634) );
  OAI222_X1 U1046 ( .A1(n38653), .A2(n35707), .B1(n38627), .B2(n35195), .C1(
        n38641), .C2(n36219), .ZN(n5640) );
  OAI222_X1 U1047 ( .A1(n37946), .A2(n35675), .B1(n37922), .B2(n35163), .C1(
        n37936), .C2(n36187), .ZN(n5641) );
  OAI222_X1 U1048 ( .A1(n38531), .A2(n35699), .B1(n38507), .B2(n35187), .C1(
        n38521), .C2(n36211), .ZN(n5642) );
  OAI222_X1 U1049 ( .A1(n37892), .A2(n35668), .B1(n37868), .B2(n35156), .C1(
        n37882), .C2(n36180), .ZN(n5590) );
  OAI222_X1 U1050 ( .A1(n38465), .A2(n35692), .B1(n38282), .B2(n35172), .C1(
        n38110), .C2(n36196), .ZN(n5591) );
  OAI222_X1 U1051 ( .A1(n38129), .A2(n35684), .B1(n38477), .B2(n35180), .C1(
        n38305), .C2(n36204), .ZN(n5592) );
  OAI222_X1 U1052 ( .A1(n38653), .A2(n35708), .B1(n38627), .B2(n35196), .C1(
        n38641), .C2(n36220), .ZN(n5598) );
  OAI222_X1 U1053 ( .A1(n37946), .A2(n35676), .B1(n37922), .B2(n35164), .C1(
        n37936), .C2(n36188), .ZN(n5599) );
  OAI222_X1 U1054 ( .A1(n38531), .A2(n35700), .B1(n38507), .B2(n35188), .C1(
        n38521), .C2(n36212), .ZN(n5600) );
  OAI222_X1 U1055 ( .A1(n37892), .A2(n35669), .B1(n37868), .B2(n35157), .C1(
        n37882), .C2(n36181), .ZN(n5527) );
  OAI222_X1 U1056 ( .A1(n38465), .A2(n35693), .B1(n38282), .B2(n35173), .C1(
        n38110), .C2(n36197), .ZN(n5530) );
  OAI222_X1 U1057 ( .A1(n38129), .A2(n35685), .B1(n38477), .B2(n35181), .C1(
        n38305), .C2(n36205), .ZN(n5533) );
  OAI222_X1 U1058 ( .A1(n38653), .A2(n35709), .B1(n38627), .B2(n35197), .C1(
        n38641), .C2(n36221), .ZN(n5539) );
  OAI222_X1 U1059 ( .A1(n37946), .A2(n35677), .B1(n37922), .B2(n35165), .C1(
        n37936), .C2(n36189), .ZN(n5541) );
  OAI222_X1 U1060 ( .A1(n38531), .A2(n35701), .B1(n38507), .B2(n35189), .C1(
        n38521), .C2(n36213), .ZN(n5542) );
  OAI222_X1 U1061 ( .A1(n37894), .A2(n35710), .B1(n37870), .B2(n35198), .C1(
        n37880), .C2(n36222), .ZN(n9576) );
  OAI222_X1 U1062 ( .A1(n38467), .A2(n35782), .B1(n38284), .B2(n35246), .C1(
        n38108), .C2(n36270), .ZN(n9582) );
  OAI222_X1 U1063 ( .A1(n38131), .A2(n35758), .B1(n38479), .B2(n35270), .C1(
        n38303), .C2(n36294), .ZN(n9588) );
  OAI222_X1 U1064 ( .A1(n38651), .A2(n35830), .B1(n38629), .B2(n35318), .C1(
        n38639), .C2(n36342), .ZN(n9598) );
  OAI222_X1 U1065 ( .A1(n37948), .A2(n35734), .B1(n37924), .B2(n35222), .C1(
        n37934), .C2(n36246), .ZN(n9600) );
  OAI222_X1 U1066 ( .A1(n38533), .A2(n35806), .B1(n38509), .B2(n35294), .C1(
        n38519), .C2(n36318), .ZN(n9606) );
  OAI222_X1 U1067 ( .A1(n37894), .A2(n35711), .B1(n37870), .B2(n35199), .C1(
        n37880), .C2(n36223), .ZN(n9528) );
  OAI222_X1 U1068 ( .A1(n38467), .A2(n35783), .B1(n38284), .B2(n35247), .C1(
        n38108), .C2(n36271), .ZN(n9529) );
  OAI222_X1 U1069 ( .A1(n38131), .A2(n35759), .B1(n38479), .B2(n35271), .C1(
        n38303), .C2(n36295), .ZN(n9530) );
  OAI222_X1 U1070 ( .A1(n38651), .A2(n35831), .B1(n38629), .B2(n35319), .C1(
        n38639), .C2(n36343), .ZN(n9536) );
  OAI222_X1 U1071 ( .A1(n37948), .A2(n35735), .B1(n37924), .B2(n35223), .C1(
        n37934), .C2(n36247), .ZN(n9537) );
  OAI222_X1 U1072 ( .A1(n38533), .A2(n35807), .B1(n38509), .B2(n35295), .C1(
        n38519), .C2(n36319), .ZN(n9538) );
  OAI222_X1 U1073 ( .A1(n37894), .A2(n35712), .B1(n37870), .B2(n35200), .C1(
        n37880), .C2(n36224), .ZN(n9486) );
  OAI222_X1 U1074 ( .A1(n38467), .A2(n35784), .B1(n38284), .B2(n35248), .C1(
        n38108), .C2(n36272), .ZN(n9487) );
  OAI222_X1 U1075 ( .A1(n38131), .A2(n35760), .B1(n38479), .B2(n35272), .C1(
        n38303), .C2(n36296), .ZN(n9488) );
  OAI222_X1 U1076 ( .A1(n38651), .A2(n35832), .B1(n38629), .B2(n35320), .C1(
        n38639), .C2(n36344), .ZN(n9494) );
  OAI222_X1 U1077 ( .A1(n37948), .A2(n35736), .B1(n37924), .B2(n35224), .C1(
        n37934), .C2(n36248), .ZN(n9495) );
  OAI222_X1 U1078 ( .A1(n38533), .A2(n35808), .B1(n38509), .B2(n35296), .C1(
        n38519), .C2(n36320), .ZN(n9496) );
  OAI222_X1 U1079 ( .A1(n37894), .A2(n35713), .B1(n37870), .B2(n35201), .C1(
        n37880), .C2(n36225), .ZN(n9444) );
  OAI222_X1 U1080 ( .A1(n38467), .A2(n35785), .B1(n38284), .B2(n35249), .C1(
        n38108), .C2(n36273), .ZN(n9445) );
  OAI222_X1 U1081 ( .A1(n38131), .A2(n35761), .B1(n38479), .B2(n35273), .C1(
        n38303), .C2(n36297), .ZN(n9446) );
  OAI222_X1 U1082 ( .A1(n38651), .A2(n35833), .B1(n38629), .B2(n35321), .C1(
        n38639), .C2(n36345), .ZN(n9452) );
  OAI222_X1 U1083 ( .A1(n37948), .A2(n35737), .B1(n37924), .B2(n35225), .C1(
        n37934), .C2(n36249), .ZN(n9453) );
  OAI222_X1 U1084 ( .A1(n38533), .A2(n35809), .B1(n38509), .B2(n35297), .C1(
        n38519), .C2(n36321), .ZN(n9454) );
  OAI222_X1 U1085 ( .A1(n37894), .A2(n35714), .B1(n37870), .B2(n35202), .C1(
        n37880), .C2(n36226), .ZN(n9402) );
  OAI222_X1 U1086 ( .A1(n38467), .A2(n35786), .B1(n38284), .B2(n35250), .C1(
        n38108), .C2(n36274), .ZN(n9403) );
  OAI222_X1 U1087 ( .A1(n38131), .A2(n35762), .B1(n38479), .B2(n35274), .C1(
        n38303), .C2(n36298), .ZN(n9404) );
  OAI222_X1 U1088 ( .A1(n38651), .A2(n35834), .B1(n38629), .B2(n35322), .C1(
        n38639), .C2(n36346), .ZN(n9410) );
  OAI222_X1 U1089 ( .A1(n37948), .A2(n35738), .B1(n37924), .B2(n35226), .C1(
        n37934), .C2(n36250), .ZN(n9411) );
  OAI222_X1 U1090 ( .A1(n38533), .A2(n35810), .B1(n38509), .B2(n35298), .C1(
        n38519), .C2(n36322), .ZN(n9412) );
  OAI222_X1 U1091 ( .A1(n37894), .A2(n35715), .B1(n37870), .B2(n35203), .C1(
        n37880), .C2(n36227), .ZN(n9360) );
  OAI222_X1 U1092 ( .A1(n38467), .A2(n35787), .B1(n38284), .B2(n35251), .C1(
        n38108), .C2(n36275), .ZN(n9361) );
  OAI222_X1 U1093 ( .A1(n38131), .A2(n35763), .B1(n38479), .B2(n35275), .C1(
        n38303), .C2(n36299), .ZN(n9362) );
  OAI222_X1 U1094 ( .A1(n38651), .A2(n35835), .B1(n38629), .B2(n35323), .C1(
        n38639), .C2(n36347), .ZN(n9368) );
  OAI222_X1 U1095 ( .A1(n37948), .A2(n35739), .B1(n37924), .B2(n35227), .C1(
        n37934), .C2(n36251), .ZN(n9369) );
  OAI222_X1 U1096 ( .A1(n38533), .A2(n35811), .B1(n38509), .B2(n35299), .C1(
        n38519), .C2(n36323), .ZN(n9370) );
  OAI222_X1 U1097 ( .A1(n37894), .A2(n35716), .B1(n37870), .B2(n35204), .C1(
        n37880), .C2(n36228), .ZN(n9318) );
  OAI222_X1 U1098 ( .A1(n38467), .A2(n35788), .B1(n38284), .B2(n35252), .C1(
        n38108), .C2(n36276), .ZN(n9319) );
  OAI222_X1 U1099 ( .A1(n38131), .A2(n35764), .B1(n38479), .B2(n35276), .C1(
        n38303), .C2(n36300), .ZN(n9320) );
  OAI222_X1 U1100 ( .A1(n38651), .A2(n35836), .B1(n38629), .B2(n35324), .C1(
        n38639), .C2(n36348), .ZN(n9326) );
  OAI222_X1 U1101 ( .A1(n37948), .A2(n35740), .B1(n37924), .B2(n35228), .C1(
        n37934), .C2(n36252), .ZN(n9327) );
  OAI222_X1 U1102 ( .A1(n38533), .A2(n35812), .B1(n38509), .B2(n35300), .C1(
        n38519), .C2(n36324), .ZN(n9328) );
  OAI222_X1 U1103 ( .A1(n37894), .A2(n35717), .B1(n37870), .B2(n35205), .C1(
        n37880), .C2(n36229), .ZN(n9276) );
  OAI222_X1 U1104 ( .A1(n38467), .A2(n35789), .B1(n38284), .B2(n35253), .C1(
        n38108), .C2(n36277), .ZN(n9277) );
  OAI222_X1 U1105 ( .A1(n38131), .A2(n35765), .B1(n38479), .B2(n35277), .C1(
        n38303), .C2(n36301), .ZN(n9278) );
  OAI222_X1 U1106 ( .A1(n38651), .A2(n35837), .B1(n38629), .B2(n35325), .C1(
        n38639), .C2(n36349), .ZN(n9284) );
  OAI222_X1 U1107 ( .A1(n37948), .A2(n35741), .B1(n37924), .B2(n35229), .C1(
        n37934), .C2(n36253), .ZN(n9285) );
  OAI222_X1 U1108 ( .A1(n38533), .A2(n35813), .B1(n38509), .B2(n35301), .C1(
        n38519), .C2(n36325), .ZN(n9286) );
  OAI222_X1 U1109 ( .A1(n37894), .A2(n35718), .B1(n37870), .B2(n35206), .C1(
        n37880), .C2(n36230), .ZN(n6642) );
  OAI222_X1 U1110 ( .A1(n38467), .A2(n35790), .B1(n38284), .B2(n35254), .C1(
        n38108), .C2(n36278), .ZN(n6643) );
  OAI222_X1 U1111 ( .A1(n38131), .A2(n35766), .B1(n38479), .B2(n35278), .C1(
        n38303), .C2(n36302), .ZN(n6644) );
  OAI222_X1 U1112 ( .A1(n38651), .A2(n35838), .B1(n38629), .B2(n35326), .C1(
        n38639), .C2(n36350), .ZN(n6650) );
  OAI222_X1 U1113 ( .A1(n37948), .A2(n35742), .B1(n37924), .B2(n35230), .C1(
        n37934), .C2(n36254), .ZN(n6651) );
  OAI222_X1 U1114 ( .A1(n38533), .A2(n35814), .B1(n38509), .B2(n35302), .C1(
        n38519), .C2(n36326), .ZN(n6652) );
  OAI222_X1 U1115 ( .A1(n37893), .A2(n35719), .B1(n37869), .B2(n35207), .C1(
        n37880), .C2(n36231), .ZN(n6600) );
  OAI222_X1 U1116 ( .A1(n38466), .A2(n35791), .B1(n38283), .B2(n35255), .C1(
        n38108), .C2(n36279), .ZN(n6601) );
  OAI222_X1 U1117 ( .A1(n38130), .A2(n35767), .B1(n38478), .B2(n35279), .C1(
        n38303), .C2(n36303), .ZN(n6602) );
  OAI222_X1 U1118 ( .A1(n38651), .A2(n35839), .B1(n38628), .B2(n35327), .C1(
        n38639), .C2(n36351), .ZN(n6608) );
  OAI222_X1 U1119 ( .A1(n37947), .A2(n35743), .B1(n37923), .B2(n35231), .C1(
        n37934), .C2(n36255), .ZN(n6609) );
  OAI222_X1 U1120 ( .A1(n38532), .A2(n35815), .B1(n38508), .B2(n35303), .C1(
        n38519), .C2(n36327), .ZN(n6610) );
  OAI222_X1 U1121 ( .A1(n37893), .A2(n35720), .B1(n37869), .B2(n35208), .C1(
        n37880), .C2(n36232), .ZN(n6558) );
  OAI222_X1 U1122 ( .A1(n38466), .A2(n35792), .B1(n38283), .B2(n35256), .C1(
        n38108), .C2(n36280), .ZN(n6559) );
  OAI222_X1 U1123 ( .A1(n38130), .A2(n35768), .B1(n38478), .B2(n35280), .C1(
        n38303), .C2(n36304), .ZN(n6560) );
  OAI222_X1 U1124 ( .A1(n38651), .A2(n35840), .B1(n38628), .B2(n35328), .C1(
        n38639), .C2(n36352), .ZN(n6566) );
  OAI222_X1 U1125 ( .A1(n37947), .A2(n35744), .B1(n37923), .B2(n35232), .C1(
        n37934), .C2(n36256), .ZN(n6567) );
  OAI222_X1 U1126 ( .A1(n38532), .A2(n35816), .B1(n38508), .B2(n35304), .C1(
        n38519), .C2(n36328), .ZN(n6568) );
  OAI222_X1 U1127 ( .A1(n37893), .A2(n35721), .B1(n37869), .B2(n35209), .C1(
        n37880), .C2(n36233), .ZN(n6516) );
  OAI222_X1 U1128 ( .A1(n38466), .A2(n35793), .B1(n38283), .B2(n35257), .C1(
        n38108), .C2(n36281), .ZN(n6517) );
  OAI222_X1 U1129 ( .A1(n38130), .A2(n35769), .B1(n38478), .B2(n35281), .C1(
        n38303), .C2(n36305), .ZN(n6518) );
  OAI222_X1 U1130 ( .A1(n38651), .A2(n35841), .B1(n38628), .B2(n35329), .C1(
        n38639), .C2(n36353), .ZN(n6524) );
  OAI222_X1 U1131 ( .A1(n37947), .A2(n35745), .B1(n37923), .B2(n35233), .C1(
        n37934), .C2(n36257), .ZN(n6525) );
  OAI222_X1 U1132 ( .A1(n38532), .A2(n35817), .B1(n38508), .B2(n35305), .C1(
        n38519), .C2(n36329), .ZN(n6526) );
  OAI222_X1 U1133 ( .A1(n37893), .A2(n35722), .B1(n37869), .B2(n35210), .C1(
        n37881), .C2(n36234), .ZN(n6346) );
  OAI222_X1 U1134 ( .A1(n38466), .A2(n35794), .B1(n38283), .B2(n35258), .C1(
        n38109), .C2(n36282), .ZN(n6347) );
  OAI222_X1 U1135 ( .A1(n38130), .A2(n35770), .B1(n38478), .B2(n35282), .C1(
        n38304), .C2(n36306), .ZN(n6348) );
  OAI222_X1 U1136 ( .A1(n38652), .A2(n35842), .B1(n38628), .B2(n35330), .C1(
        n38640), .C2(n36354), .ZN(n6354) );
  OAI222_X1 U1137 ( .A1(n37947), .A2(n35746), .B1(n37923), .B2(n35234), .C1(
        n37935), .C2(n36258), .ZN(n6355) );
  OAI222_X1 U1138 ( .A1(n38532), .A2(n35818), .B1(n38508), .B2(n35306), .C1(
        n38520), .C2(n36330), .ZN(n6356) );
  OAI222_X1 U1139 ( .A1(n37893), .A2(n35723), .B1(n37869), .B2(n35211), .C1(
        n37881), .C2(n36235), .ZN(n6304) );
  OAI222_X1 U1140 ( .A1(n38466), .A2(n35795), .B1(n38283), .B2(n35259), .C1(
        n38109), .C2(n36283), .ZN(n6305) );
  OAI222_X1 U1141 ( .A1(n38130), .A2(n35771), .B1(n38478), .B2(n35283), .C1(
        n38304), .C2(n36307), .ZN(n6306) );
  OAI222_X1 U1142 ( .A1(n38652), .A2(n35843), .B1(n38628), .B2(n35331), .C1(
        n38640), .C2(n36355), .ZN(n6312) );
  OAI222_X1 U1143 ( .A1(n37947), .A2(n35747), .B1(n37923), .B2(n35235), .C1(
        n37935), .C2(n36259), .ZN(n6313) );
  OAI222_X1 U1144 ( .A1(n38532), .A2(n35819), .B1(n38508), .B2(n35307), .C1(
        n38520), .C2(n36331), .ZN(n6314) );
  OAI222_X1 U1145 ( .A1(n37893), .A2(n35724), .B1(n37869), .B2(n35212), .C1(
        n37881), .C2(n36236), .ZN(n6262) );
  OAI222_X1 U1146 ( .A1(n38466), .A2(n35796), .B1(n38283), .B2(n35260), .C1(
        n38109), .C2(n36284), .ZN(n6263) );
  OAI222_X1 U1147 ( .A1(n38130), .A2(n35772), .B1(n38478), .B2(n35284), .C1(
        n38304), .C2(n36308), .ZN(n6264) );
  OAI222_X1 U1148 ( .A1(n38652), .A2(n35844), .B1(n38628), .B2(n35332), .C1(
        n38640), .C2(n36356), .ZN(n6270) );
  OAI222_X1 U1149 ( .A1(n37947), .A2(n35748), .B1(n37923), .B2(n35236), .C1(
        n37935), .C2(n36260), .ZN(n6271) );
  OAI222_X1 U1150 ( .A1(n38532), .A2(n35820), .B1(n38508), .B2(n35308), .C1(
        n38520), .C2(n36332), .ZN(n6272) );
  OAI222_X1 U1151 ( .A1(n37893), .A2(n35725), .B1(n37869), .B2(n35213), .C1(
        n37881), .C2(n36237), .ZN(n6220) );
  OAI222_X1 U1152 ( .A1(n38466), .A2(n35797), .B1(n38283), .B2(n35261), .C1(
        n38109), .C2(n36285), .ZN(n6221) );
  OAI222_X1 U1153 ( .A1(n38130), .A2(n35773), .B1(n38478), .B2(n35285), .C1(
        n38304), .C2(n36309), .ZN(n6222) );
  OAI222_X1 U1154 ( .A1(n38652), .A2(n35845), .B1(n38628), .B2(n35333), .C1(
        n38640), .C2(n36357), .ZN(n6228) );
  OAI222_X1 U1155 ( .A1(n37947), .A2(n35749), .B1(n37923), .B2(n35237), .C1(
        n37935), .C2(n36261), .ZN(n6229) );
  OAI222_X1 U1156 ( .A1(n38532), .A2(n35821), .B1(n38508), .B2(n35309), .C1(
        n38520), .C2(n36333), .ZN(n6230) );
  OAI222_X1 U1157 ( .A1(n37893), .A2(n35726), .B1(n37869), .B2(n35214), .C1(
        n37881), .C2(n36238), .ZN(n6178) );
  OAI222_X1 U1158 ( .A1(n38466), .A2(n35798), .B1(n38283), .B2(n35262), .C1(
        n38109), .C2(n36286), .ZN(n6179) );
  OAI222_X1 U1159 ( .A1(n38130), .A2(n35774), .B1(n38478), .B2(n35286), .C1(
        n38304), .C2(n36310), .ZN(n6180) );
  OAI222_X1 U1160 ( .A1(n38652), .A2(n35846), .B1(n38628), .B2(n35334), .C1(
        n38640), .C2(n36358), .ZN(n6186) );
  OAI222_X1 U1161 ( .A1(n37947), .A2(n35750), .B1(n37923), .B2(n35238), .C1(
        n37935), .C2(n36262), .ZN(n6187) );
  OAI222_X1 U1162 ( .A1(n38532), .A2(n35822), .B1(n38508), .B2(n35310), .C1(
        n38520), .C2(n36334), .ZN(n6188) );
  OAI222_X1 U1163 ( .A1(n37893), .A2(n35727), .B1(n37869), .B2(n35215), .C1(
        n37881), .C2(n36239), .ZN(n6136) );
  OAI222_X1 U1164 ( .A1(n38466), .A2(n35799), .B1(n38283), .B2(n35263), .C1(
        n38109), .C2(n36287), .ZN(n6137) );
  OAI222_X1 U1165 ( .A1(n38130), .A2(n35775), .B1(n38478), .B2(n35287), .C1(
        n38304), .C2(n36311), .ZN(n6138) );
  OAI222_X1 U1166 ( .A1(n38652), .A2(n35847), .B1(n38628), .B2(n35335), .C1(
        n38640), .C2(n36359), .ZN(n6144) );
  OAI222_X1 U1167 ( .A1(n37947), .A2(n35751), .B1(n37923), .B2(n35239), .C1(
        n37935), .C2(n36263), .ZN(n6145) );
  OAI222_X1 U1168 ( .A1(n38532), .A2(n35823), .B1(n38508), .B2(n35311), .C1(
        n38520), .C2(n36335), .ZN(n6146) );
  OAI222_X1 U1169 ( .A1(n37893), .A2(n35728), .B1(n37869), .B2(n35216), .C1(
        n37881), .C2(n36240), .ZN(n6094) );
  OAI222_X1 U1170 ( .A1(n38466), .A2(n35800), .B1(n38283), .B2(n35264), .C1(
        n38109), .C2(n36288), .ZN(n6095) );
  OAI222_X1 U1171 ( .A1(n38130), .A2(n35776), .B1(n38478), .B2(n35288), .C1(
        n38304), .C2(n36312), .ZN(n6096) );
  OAI222_X1 U1172 ( .A1(n38652), .A2(n35848), .B1(n38628), .B2(n35336), .C1(
        n38640), .C2(n36360), .ZN(n6102) );
  OAI222_X1 U1173 ( .A1(n37947), .A2(n35752), .B1(n37923), .B2(n35240), .C1(
        n37935), .C2(n36264), .ZN(n6103) );
  OAI222_X1 U1174 ( .A1(n38532), .A2(n35824), .B1(n38508), .B2(n35312), .C1(
        n38520), .C2(n36336), .ZN(n6104) );
  OAI222_X1 U1175 ( .A1(n37893), .A2(n35729), .B1(n37869), .B2(n35217), .C1(
        n37881), .C2(n36241), .ZN(n6052) );
  OAI222_X1 U1176 ( .A1(n38466), .A2(n35801), .B1(n38283), .B2(n35265), .C1(
        n38109), .C2(n36289), .ZN(n6053) );
  OAI222_X1 U1177 ( .A1(n38130), .A2(n35777), .B1(n38478), .B2(n35289), .C1(
        n38304), .C2(n36313), .ZN(n6054) );
  OAI222_X1 U1178 ( .A1(n38652), .A2(n35849), .B1(n38628), .B2(n35337), .C1(
        n38640), .C2(n36361), .ZN(n6060) );
  OAI222_X1 U1179 ( .A1(n37947), .A2(n35753), .B1(n37923), .B2(n35241), .C1(
        n37935), .C2(n36265), .ZN(n6061) );
  OAI222_X1 U1180 ( .A1(n38532), .A2(n35825), .B1(n38508), .B2(n35313), .C1(
        n38520), .C2(n36337), .ZN(n6062) );
  OAI222_X1 U1181 ( .A1(n37893), .A2(n35730), .B1(n37869), .B2(n35218), .C1(
        n37881), .C2(n36242), .ZN(n6010) );
  OAI222_X1 U1182 ( .A1(n38466), .A2(n35802), .B1(n38283), .B2(n35266), .C1(
        n38109), .C2(n36290), .ZN(n6011) );
  OAI222_X1 U1183 ( .A1(n38130), .A2(n35778), .B1(n38478), .B2(n35290), .C1(
        n38304), .C2(n36314), .ZN(n6012) );
  OAI222_X1 U1184 ( .A1(n38652), .A2(n35850), .B1(n38628), .B2(n35338), .C1(
        n38640), .C2(n36362), .ZN(n6018) );
  OAI222_X1 U1185 ( .A1(n37947), .A2(n35754), .B1(n37923), .B2(n35242), .C1(
        n37935), .C2(n36266), .ZN(n6019) );
  OAI222_X1 U1186 ( .A1(n38532), .A2(n35826), .B1(n38508), .B2(n35314), .C1(
        n38520), .C2(n36338), .ZN(n6020) );
  OAI222_X1 U1187 ( .A1(n37892), .A2(n35731), .B1(n37868), .B2(n35219), .C1(
        n37881), .C2(n36243), .ZN(n5968) );
  OAI222_X1 U1188 ( .A1(n38465), .A2(n35803), .B1(n38282), .B2(n35267), .C1(
        n38109), .C2(n36291), .ZN(n5969) );
  OAI222_X1 U1189 ( .A1(n38129), .A2(n35779), .B1(n38477), .B2(n35291), .C1(
        n38304), .C2(n36315), .ZN(n5970) );
  OAI222_X1 U1190 ( .A1(n38652), .A2(n35851), .B1(n38627), .B2(n35339), .C1(
        n38640), .C2(n36363), .ZN(n5976) );
  OAI222_X1 U1191 ( .A1(n37946), .A2(n35755), .B1(n37922), .B2(n35243), .C1(
        n37935), .C2(n36267), .ZN(n5977) );
  OAI222_X1 U1192 ( .A1(n38531), .A2(n35827), .B1(n38507), .B2(n35315), .C1(
        n38520), .C2(n36339), .ZN(n5978) );
  OAI222_X1 U1193 ( .A1(n37892), .A2(n35732), .B1(n37868), .B2(n35220), .C1(
        n37881), .C2(n36244), .ZN(n5926) );
  OAI222_X1 U1194 ( .A1(n38465), .A2(n35804), .B1(n38282), .B2(n35268), .C1(
        n38109), .C2(n36292), .ZN(n5927) );
  OAI222_X1 U1195 ( .A1(n38129), .A2(n35780), .B1(n38477), .B2(n35292), .C1(
        n38304), .C2(n36316), .ZN(n5928) );
  OAI222_X1 U1196 ( .A1(n38652), .A2(n35852), .B1(n38627), .B2(n35340), .C1(
        n38640), .C2(n36364), .ZN(n5934) );
  OAI222_X1 U1197 ( .A1(n37946), .A2(n35756), .B1(n37922), .B2(n35244), .C1(
        n37935), .C2(n36268), .ZN(n5935) );
  OAI222_X1 U1198 ( .A1(n38531), .A2(n35828), .B1(n38507), .B2(n35316), .C1(
        n38520), .C2(n36340), .ZN(n5936) );
  OAI222_X1 U1199 ( .A1(n37892), .A2(n35733), .B1(n37868), .B2(n35221), .C1(
        n37881), .C2(n36245), .ZN(n5884) );
  OAI222_X1 U1200 ( .A1(n38465), .A2(n35805), .B1(n38282), .B2(n35269), .C1(
        n38109), .C2(n36293), .ZN(n5885) );
  OAI222_X1 U1201 ( .A1(n38129), .A2(n35781), .B1(n38477), .B2(n35293), .C1(
        n38304), .C2(n36317), .ZN(n5886) );
  OAI222_X1 U1202 ( .A1(n38652), .A2(n35853), .B1(n38627), .B2(n35341), .C1(
        n38640), .C2(n36365), .ZN(n5892) );
  OAI222_X1 U1203 ( .A1(n37946), .A2(n35757), .B1(n37922), .B2(n35245), .C1(
        n37935), .C2(n36269), .ZN(n5893) );
  OAI222_X1 U1204 ( .A1(n38531), .A2(n35829), .B1(n38507), .B2(n35317), .C1(
        n38520), .C2(n36341), .ZN(n5894) );
  OAI21_X1 U1205 ( .B1(n5016), .B2(n9560), .A(n38919), .ZN(n5508) );
  BUF_X1 U1206 ( .A(n2739), .Z(n38683) );
  BUF_X1 U1207 ( .A(n2737), .Z(n38690) );
  BUF_X1 U1208 ( .A(n2735), .Z(n38697) );
  BUF_X1 U1209 ( .A(n2733), .Z(n38704) );
  BUF_X1 U1210 ( .A(n2731), .Z(n38711) );
  BUF_X1 U1211 ( .A(n2729), .Z(n38718) );
  BUF_X1 U1212 ( .A(n2727), .Z(n38725) );
  BUF_X1 U1213 ( .A(n2725), .Z(n38732) );
  BUF_X1 U1214 ( .A(n2723), .Z(n38739) );
  BUF_X1 U1215 ( .A(n2721), .Z(n38746) );
  BUF_X1 U1216 ( .A(n2719), .Z(n38753) );
  BUF_X1 U1217 ( .A(n2717), .Z(n38760) );
  BUF_X1 U1218 ( .A(n2739), .Z(n38682) );
  BUF_X1 U1219 ( .A(n2737), .Z(n38689) );
  BUF_X1 U1220 ( .A(n2735), .Z(n38696) );
  BUF_X1 U1221 ( .A(n2733), .Z(n38703) );
  BUF_X1 U1222 ( .A(n2731), .Z(n38710) );
  BUF_X1 U1223 ( .A(n2729), .Z(n38717) );
  BUF_X1 U1224 ( .A(n2727), .Z(n38724) );
  BUF_X1 U1225 ( .A(n2725), .Z(n38731) );
  BUF_X1 U1226 ( .A(n2723), .Z(n38738) );
  BUF_X1 U1227 ( .A(n2721), .Z(n38745) );
  BUF_X1 U1228 ( .A(n2719), .Z(n38752) );
  BUF_X1 U1229 ( .A(n2717), .Z(n38759) );
  BUF_X1 U1230 ( .A(n2739), .Z(n38681) );
  BUF_X1 U1231 ( .A(n2737), .Z(n38688) );
  BUF_X1 U1232 ( .A(n2735), .Z(n38695) );
  BUF_X1 U1233 ( .A(n2733), .Z(n38702) );
  BUF_X1 U1234 ( .A(n2731), .Z(n38709) );
  BUF_X1 U1235 ( .A(n2729), .Z(n38716) );
  BUF_X1 U1236 ( .A(n2727), .Z(n38723) );
  BUF_X1 U1237 ( .A(n2725), .Z(n38730) );
  BUF_X1 U1238 ( .A(n2723), .Z(n38737) );
  BUF_X1 U1239 ( .A(n2721), .Z(n38744) );
  BUF_X1 U1240 ( .A(n2719), .Z(n38751) );
  BUF_X1 U1241 ( .A(n2717), .Z(n38758) );
  BUF_X1 U1242 ( .A(n2739), .Z(n38680) );
  BUF_X1 U1243 ( .A(n2737), .Z(n38687) );
  BUF_X1 U1244 ( .A(n2735), .Z(n38694) );
  BUF_X1 U1245 ( .A(n2733), .Z(n38701) );
  BUF_X1 U1246 ( .A(n2731), .Z(n38708) );
  BUF_X1 U1247 ( .A(n2729), .Z(n38715) );
  BUF_X1 U1248 ( .A(n2727), .Z(n38722) );
  BUF_X1 U1249 ( .A(n2725), .Z(n38729) );
  BUF_X1 U1250 ( .A(n2723), .Z(n38736) );
  BUF_X1 U1251 ( .A(n2721), .Z(n38743) );
  BUF_X1 U1252 ( .A(n2719), .Z(n38750) );
  BUF_X1 U1253 ( .A(n2717), .Z(n38757) );
  BUF_X1 U1254 ( .A(n2739), .Z(n38679) );
  BUF_X1 U1255 ( .A(n2737), .Z(n38686) );
  BUF_X1 U1256 ( .A(n2735), .Z(n38693) );
  BUF_X1 U1257 ( .A(n2733), .Z(n38700) );
  BUF_X1 U1258 ( .A(n2731), .Z(n38707) );
  BUF_X1 U1259 ( .A(n2729), .Z(n38714) );
  BUF_X1 U1260 ( .A(n2727), .Z(n38721) );
  BUF_X1 U1261 ( .A(n2725), .Z(n38728) );
  BUF_X1 U1262 ( .A(n2723), .Z(n38735) );
  BUF_X1 U1263 ( .A(n2721), .Z(n38742) );
  BUF_X1 U1264 ( .A(n2719), .Z(n38749) );
  BUF_X1 U1265 ( .A(n2717), .Z(n38756) );
  BUF_X1 U1266 ( .A(n2739), .Z(n38678) );
  BUF_X1 U1267 ( .A(n2737), .Z(n38685) );
  BUF_X1 U1268 ( .A(n2735), .Z(n38692) );
  BUF_X1 U1269 ( .A(n2733), .Z(n38699) );
  BUF_X1 U1270 ( .A(n2731), .Z(n38706) );
  BUF_X1 U1271 ( .A(n2729), .Z(n38713) );
  BUF_X1 U1272 ( .A(n2727), .Z(n38720) );
  BUF_X1 U1273 ( .A(n2725), .Z(n38727) );
  BUF_X1 U1274 ( .A(n2723), .Z(n38734) );
  BUF_X1 U1275 ( .A(n2721), .Z(n38741) );
  BUF_X1 U1276 ( .A(n2719), .Z(n38748) );
  BUF_X1 U1277 ( .A(n2717), .Z(n38755) );
  BUF_X1 U1278 ( .A(n2715), .Z(n38767) );
  BUF_X1 U1279 ( .A(n2713), .Z(n38774) );
  BUF_X1 U1280 ( .A(n2711), .Z(n38781) );
  BUF_X1 U1281 ( .A(n2709), .Z(n38788) );
  BUF_X1 U1282 ( .A(n2707), .Z(n38795) );
  BUF_X1 U1283 ( .A(n2705), .Z(n38802) );
  BUF_X1 U1284 ( .A(n2703), .Z(n38809) );
  BUF_X1 U1285 ( .A(n2701), .Z(n38816) );
  BUF_X1 U1286 ( .A(n2699), .Z(n38823) );
  BUF_X1 U1287 ( .A(n2697), .Z(n38830) );
  BUF_X1 U1288 ( .A(n2695), .Z(n38837) );
  BUF_X1 U1289 ( .A(n2693), .Z(n38844) );
  BUF_X1 U1290 ( .A(n2691), .Z(n38851) );
  BUF_X1 U1291 ( .A(n2689), .Z(n38858) );
  BUF_X1 U1292 ( .A(n2687), .Z(n38865) );
  BUF_X1 U1293 ( .A(n2685), .Z(n38872) );
  BUF_X1 U1294 ( .A(n2683), .Z(n38879) );
  BUF_X1 U1295 ( .A(n2681), .Z(n38886) );
  BUF_X1 U1296 ( .A(n2679), .Z(n38893) );
  BUF_X1 U1297 ( .A(n2677), .Z(n38900) );
  BUF_X1 U1298 ( .A(n2715), .Z(n38766) );
  BUF_X1 U1299 ( .A(n2713), .Z(n38773) );
  BUF_X1 U1300 ( .A(n2711), .Z(n38780) );
  BUF_X1 U1301 ( .A(n2709), .Z(n38787) );
  BUF_X1 U1302 ( .A(n2707), .Z(n38794) );
  BUF_X1 U1303 ( .A(n2705), .Z(n38801) );
  BUF_X1 U1304 ( .A(n2703), .Z(n38808) );
  BUF_X1 U1305 ( .A(n2701), .Z(n38815) );
  BUF_X1 U1306 ( .A(n2699), .Z(n38822) );
  BUF_X1 U1307 ( .A(n2697), .Z(n38829) );
  BUF_X1 U1308 ( .A(n2695), .Z(n38836) );
  BUF_X1 U1309 ( .A(n2693), .Z(n38843) );
  BUF_X1 U1310 ( .A(n2691), .Z(n38850) );
  BUF_X1 U1311 ( .A(n2689), .Z(n38857) );
  BUF_X1 U1312 ( .A(n2687), .Z(n38864) );
  BUF_X1 U1313 ( .A(n2685), .Z(n38871) );
  BUF_X1 U1314 ( .A(n2683), .Z(n38878) );
  BUF_X1 U1315 ( .A(n2681), .Z(n38885) );
  BUF_X1 U1316 ( .A(n2679), .Z(n38892) );
  BUF_X1 U1317 ( .A(n2677), .Z(n38899) );
  BUF_X1 U1318 ( .A(n2715), .Z(n38765) );
  BUF_X1 U1319 ( .A(n2713), .Z(n38772) );
  BUF_X1 U1320 ( .A(n2711), .Z(n38779) );
  BUF_X1 U1321 ( .A(n2709), .Z(n38786) );
  BUF_X1 U1322 ( .A(n2707), .Z(n38793) );
  BUF_X1 U1323 ( .A(n2705), .Z(n38800) );
  BUF_X1 U1324 ( .A(n2703), .Z(n38807) );
  BUF_X1 U1325 ( .A(n2701), .Z(n38814) );
  BUF_X1 U1326 ( .A(n2699), .Z(n38821) );
  BUF_X1 U1327 ( .A(n2697), .Z(n38828) );
  BUF_X1 U1328 ( .A(n2695), .Z(n38835) );
  BUF_X1 U1329 ( .A(n2693), .Z(n38842) );
  BUF_X1 U1330 ( .A(n2691), .Z(n38849) );
  BUF_X1 U1331 ( .A(n2689), .Z(n38856) );
  BUF_X1 U1332 ( .A(n2687), .Z(n38863) );
  BUF_X1 U1333 ( .A(n2685), .Z(n38870) );
  BUF_X1 U1334 ( .A(n2683), .Z(n38877) );
  BUF_X1 U1335 ( .A(n2681), .Z(n38884) );
  BUF_X1 U1336 ( .A(n2679), .Z(n38891) );
  BUF_X1 U1337 ( .A(n2677), .Z(n38898) );
  BUF_X1 U1338 ( .A(n2715), .Z(n38764) );
  BUF_X1 U1339 ( .A(n2713), .Z(n38771) );
  BUF_X1 U1340 ( .A(n2711), .Z(n38778) );
  BUF_X1 U1341 ( .A(n2709), .Z(n38785) );
  BUF_X1 U1342 ( .A(n2707), .Z(n38792) );
  BUF_X1 U1343 ( .A(n2705), .Z(n38799) );
  BUF_X1 U1344 ( .A(n2703), .Z(n38806) );
  BUF_X1 U1345 ( .A(n2701), .Z(n38813) );
  BUF_X1 U1346 ( .A(n2699), .Z(n38820) );
  BUF_X1 U1347 ( .A(n2697), .Z(n38827) );
  BUF_X1 U1348 ( .A(n2695), .Z(n38834) );
  BUF_X1 U1349 ( .A(n2693), .Z(n38841) );
  BUF_X1 U1350 ( .A(n2691), .Z(n38848) );
  BUF_X1 U1351 ( .A(n2689), .Z(n38855) );
  BUF_X1 U1352 ( .A(n2687), .Z(n38862) );
  BUF_X1 U1353 ( .A(n2685), .Z(n38869) );
  BUF_X1 U1354 ( .A(n2683), .Z(n38876) );
  BUF_X1 U1355 ( .A(n2681), .Z(n38883) );
  BUF_X1 U1356 ( .A(n2679), .Z(n38890) );
  BUF_X1 U1357 ( .A(n2677), .Z(n38897) );
  BUF_X1 U1358 ( .A(n2715), .Z(n38763) );
  BUF_X1 U1359 ( .A(n2713), .Z(n38770) );
  BUF_X1 U1360 ( .A(n2711), .Z(n38777) );
  BUF_X1 U1361 ( .A(n2709), .Z(n38784) );
  BUF_X1 U1362 ( .A(n2707), .Z(n38791) );
  BUF_X1 U1363 ( .A(n2705), .Z(n38798) );
  BUF_X1 U1364 ( .A(n2703), .Z(n38805) );
  BUF_X1 U1365 ( .A(n2701), .Z(n38812) );
  BUF_X1 U1366 ( .A(n2699), .Z(n38819) );
  BUF_X1 U1367 ( .A(n2697), .Z(n38826) );
  BUF_X1 U1368 ( .A(n2695), .Z(n38833) );
  BUF_X1 U1369 ( .A(n2693), .Z(n38840) );
  BUF_X1 U1370 ( .A(n2691), .Z(n38847) );
  BUF_X1 U1371 ( .A(n2689), .Z(n38854) );
  BUF_X1 U1372 ( .A(n2687), .Z(n38861) );
  BUF_X1 U1373 ( .A(n2685), .Z(n38868) );
  BUF_X1 U1374 ( .A(n2683), .Z(n38875) );
  BUF_X1 U1375 ( .A(n2681), .Z(n38882) );
  BUF_X1 U1376 ( .A(n2679), .Z(n38889) );
  BUF_X1 U1377 ( .A(n2677), .Z(n38896) );
  BUF_X1 U1378 ( .A(n2715), .Z(n38762) );
  BUF_X1 U1379 ( .A(n2713), .Z(n38769) );
  BUF_X1 U1380 ( .A(n2711), .Z(n38776) );
  BUF_X1 U1381 ( .A(n2709), .Z(n38783) );
  BUF_X1 U1382 ( .A(n2707), .Z(n38790) );
  BUF_X1 U1383 ( .A(n2705), .Z(n38797) );
  BUF_X1 U1384 ( .A(n2703), .Z(n38804) );
  BUF_X1 U1385 ( .A(n2701), .Z(n38811) );
  BUF_X1 U1386 ( .A(n2699), .Z(n38818) );
  BUF_X1 U1387 ( .A(n2697), .Z(n38825) );
  BUF_X1 U1388 ( .A(n2695), .Z(n38832) );
  BUF_X1 U1389 ( .A(n2693), .Z(n38839) );
  BUF_X1 U1390 ( .A(n2691), .Z(n38846) );
  BUF_X1 U1391 ( .A(n2689), .Z(n38853) );
  BUF_X1 U1392 ( .A(n2687), .Z(n38860) );
  BUF_X1 U1393 ( .A(n2685), .Z(n38867) );
  BUF_X1 U1394 ( .A(n2683), .Z(n38874) );
  BUF_X1 U1395 ( .A(n2681), .Z(n38881) );
  BUF_X1 U1396 ( .A(n2679), .Z(n38888) );
  BUF_X1 U1397 ( .A(n2677), .Z(n38895) );
  NAND2_X1 U1398 ( .A1(n38918), .A2(n2812), .ZN(n2741) );
  OAI22_X1 U1399 ( .A1(n37822), .A2(n38851), .B1(n5439), .B2(n35342), .ZN(
        n6795) );
  OAI22_X1 U1400 ( .A1(n37823), .A2(n38858), .B1(n5439), .B2(n35351), .ZN(
        n6796) );
  OAI22_X1 U1401 ( .A1(n37823), .A2(n38865), .B1(n5439), .B2(n35360), .ZN(
        n6797) );
  OAI22_X1 U1402 ( .A1(n37823), .A2(n38872), .B1(n37817), .B2(n35369), .ZN(
        n6798) );
  OAI22_X1 U1403 ( .A1(n37823), .A2(n38879), .B1(n37817), .B2(n35378), .ZN(
        n6799) );
  OAI22_X1 U1404 ( .A1(n37823), .A2(n38886), .B1(n37817), .B2(n35387), .ZN(
        n6800) );
  OAI22_X1 U1405 ( .A1(n37824), .A2(n38893), .B1(n37817), .B2(n35396), .ZN(
        n6801) );
  OAI22_X1 U1406 ( .A1(n37824), .A2(n38900), .B1(n5439), .B2(n35405), .ZN(
        n6802) );
  OAI22_X1 U1407 ( .A1(n37834), .A2(n38851), .B1(n5404), .B2(n36366), .ZN(
        n6827) );
  OAI22_X1 U1408 ( .A1(n37835), .A2(n38858), .B1(n5404), .B2(n36375), .ZN(
        n6828) );
  OAI22_X1 U1409 ( .A1(n37835), .A2(n38865), .B1(n5404), .B2(n36384), .ZN(
        n6829) );
  OAI22_X1 U1410 ( .A1(n37835), .A2(n38872), .B1(n37829), .B2(n36393), .ZN(
        n6830) );
  OAI22_X1 U1411 ( .A1(n37835), .A2(n38879), .B1(n37829), .B2(n36402), .ZN(
        n6831) );
  OAI22_X1 U1412 ( .A1(n37835), .A2(n38886), .B1(n37829), .B2(n36411), .ZN(
        n6832) );
  OAI22_X1 U1413 ( .A1(n37836), .A2(n38893), .B1(n37829), .B2(n36420), .ZN(
        n6833) );
  OAI22_X1 U1414 ( .A1(n37836), .A2(n38900), .B1(n5404), .B2(n36429), .ZN(
        n6834) );
  OAI22_X1 U1415 ( .A1(n37846), .A2(n38851), .B1(n5369), .B2(n35854), .ZN(
        n6859) );
  OAI22_X1 U1416 ( .A1(n37847), .A2(n38858), .B1(n5369), .B2(n35863), .ZN(
        n6860) );
  OAI22_X1 U1417 ( .A1(n37847), .A2(n38865), .B1(n5369), .B2(n35872), .ZN(
        n6861) );
  OAI22_X1 U1418 ( .A1(n37847), .A2(n38872), .B1(n37841), .B2(n35881), .ZN(
        n6862) );
  OAI22_X1 U1419 ( .A1(n37847), .A2(n38879), .B1(n37841), .B2(n35890), .ZN(
        n6863) );
  OAI22_X1 U1420 ( .A1(n37847), .A2(n38886), .B1(n37841), .B2(n35899), .ZN(
        n6864) );
  OAI22_X1 U1421 ( .A1(n37848), .A2(n38893), .B1(n37841), .B2(n35908), .ZN(
        n6865) );
  OAI22_X1 U1422 ( .A1(n37848), .A2(n38900), .B1(n5369), .B2(n35917), .ZN(
        n6866) );
  OAI22_X1 U1423 ( .A1(n37876), .A2(n38851), .B1(n5264), .B2(n35150), .ZN(
        n6955) );
  OAI22_X1 U1424 ( .A1(n37877), .A2(n38858), .B1(n5264), .B2(n35151), .ZN(
        n6956) );
  OAI22_X1 U1425 ( .A1(n37877), .A2(n38865), .B1(n5264), .B2(n35152), .ZN(
        n6957) );
  OAI22_X1 U1426 ( .A1(n37877), .A2(n38872), .B1(n37871), .B2(n35153), .ZN(
        n6958) );
  OAI22_X1 U1427 ( .A1(n37877), .A2(n38879), .B1(n37871), .B2(n35154), .ZN(
        n6959) );
  OAI22_X1 U1428 ( .A1(n37877), .A2(n38886), .B1(n37871), .B2(n35155), .ZN(
        n6960) );
  OAI22_X1 U1429 ( .A1(n37878), .A2(n38893), .B1(n37871), .B2(n35156), .ZN(
        n6961) );
  OAI22_X1 U1430 ( .A1(n37878), .A2(n38900), .B1(n5264), .B2(n35157), .ZN(
        n6962) );
  OAI22_X1 U1431 ( .A1(n37888), .A2(n38851), .B1(n5229), .B2(n36174), .ZN(
        n6987) );
  OAI22_X1 U1432 ( .A1(n37889), .A2(n38858), .B1(n5229), .B2(n36175), .ZN(
        n6988) );
  OAI22_X1 U1433 ( .A1(n37889), .A2(n38865), .B1(n5229), .B2(n36176), .ZN(
        n6989) );
  OAI22_X1 U1434 ( .A1(n37889), .A2(n38872), .B1(n37883), .B2(n36177), .ZN(
        n6990) );
  OAI22_X1 U1435 ( .A1(n37889), .A2(n38879), .B1(n37883), .B2(n36178), .ZN(
        n6991) );
  OAI22_X1 U1436 ( .A1(n37889), .A2(n38886), .B1(n37883), .B2(n36179), .ZN(
        n6992) );
  OAI22_X1 U1437 ( .A1(n37890), .A2(n38893), .B1(n37883), .B2(n36180), .ZN(
        n6993) );
  OAI22_X1 U1438 ( .A1(n37890), .A2(n38900), .B1(n5229), .B2(n36181), .ZN(
        n6994) );
  OAI22_X1 U1439 ( .A1(n37900), .A2(n38851), .B1(n5194), .B2(n35662), .ZN(
        n7019) );
  OAI22_X1 U1440 ( .A1(n37901), .A2(n38858), .B1(n5194), .B2(n35663), .ZN(
        n7020) );
  OAI22_X1 U1441 ( .A1(n37901), .A2(n38865), .B1(n5194), .B2(n35664), .ZN(
        n7021) );
  OAI22_X1 U1442 ( .A1(n37901), .A2(n38872), .B1(n37895), .B2(n35665), .ZN(
        n7022) );
  OAI22_X1 U1443 ( .A1(n37901), .A2(n38879), .B1(n37895), .B2(n35666), .ZN(
        n7023) );
  OAI22_X1 U1444 ( .A1(n37901), .A2(n38886), .B1(n37895), .B2(n35667), .ZN(
        n7024) );
  OAI22_X1 U1445 ( .A1(n37902), .A2(n38893), .B1(n37895), .B2(n35668), .ZN(
        n7025) );
  OAI22_X1 U1446 ( .A1(n37902), .A2(n38900), .B1(n5194), .B2(n35669), .ZN(
        n7026) );
  OAI22_X1 U1447 ( .A1(n37930), .A2(n38851), .B1(n5089), .B2(n35158), .ZN(
        n7115) );
  OAI22_X1 U1448 ( .A1(n37931), .A2(n38858), .B1(n5089), .B2(n35159), .ZN(
        n7116) );
  OAI22_X1 U1449 ( .A1(n37931), .A2(n38865), .B1(n5089), .B2(n35160), .ZN(
        n7117) );
  OAI22_X1 U1450 ( .A1(n37931), .A2(n38872), .B1(n37925), .B2(n35161), .ZN(
        n7118) );
  OAI22_X1 U1451 ( .A1(n37931), .A2(n38879), .B1(n37925), .B2(n35162), .ZN(
        n7119) );
  OAI22_X1 U1452 ( .A1(n37931), .A2(n38886), .B1(n37925), .B2(n35163), .ZN(
        n7120) );
  OAI22_X1 U1453 ( .A1(n37932), .A2(n38893), .B1(n37925), .B2(n35164), .ZN(
        n7121) );
  OAI22_X1 U1454 ( .A1(n37932), .A2(n38900), .B1(n5089), .B2(n35165), .ZN(
        n7122) );
  OAI22_X1 U1455 ( .A1(n37942), .A2(n38850), .B1(n5054), .B2(n36182), .ZN(
        n7147) );
  OAI22_X1 U1456 ( .A1(n37943), .A2(n38857), .B1(n5054), .B2(n36183), .ZN(
        n7148) );
  OAI22_X1 U1457 ( .A1(n37943), .A2(n38864), .B1(n5054), .B2(n36184), .ZN(
        n7149) );
  OAI22_X1 U1458 ( .A1(n37943), .A2(n38871), .B1(n37937), .B2(n36185), .ZN(
        n7150) );
  OAI22_X1 U1459 ( .A1(n37943), .A2(n38878), .B1(n37937), .B2(n36186), .ZN(
        n7151) );
  OAI22_X1 U1460 ( .A1(n37943), .A2(n38885), .B1(n37937), .B2(n36187), .ZN(
        n7152) );
  OAI22_X1 U1461 ( .A1(n37944), .A2(n38892), .B1(n37937), .B2(n36188), .ZN(
        n7153) );
  OAI22_X1 U1462 ( .A1(n37944), .A2(n38899), .B1(n5054), .B2(n36189), .ZN(
        n7154) );
  OAI22_X1 U1463 ( .A1(n37954), .A2(n38850), .B1(n5019), .B2(n35670), .ZN(
        n7179) );
  OAI22_X1 U1464 ( .A1(n37955), .A2(n38857), .B1(n5019), .B2(n35671), .ZN(
        n7180) );
  OAI22_X1 U1465 ( .A1(n37955), .A2(n38864), .B1(n5019), .B2(n35672), .ZN(
        n7181) );
  OAI22_X1 U1466 ( .A1(n37955), .A2(n38871), .B1(n37949), .B2(n35673), .ZN(
        n7182) );
  OAI22_X1 U1467 ( .A1(n37955), .A2(n38878), .B1(n37949), .B2(n35674), .ZN(
        n7183) );
  OAI22_X1 U1468 ( .A1(n37955), .A2(n38885), .B1(n37949), .B2(n35675), .ZN(
        n7184) );
  OAI22_X1 U1469 ( .A1(n37956), .A2(n38892), .B1(n37949), .B2(n35676), .ZN(
        n7185) );
  OAI22_X1 U1470 ( .A1(n37956), .A2(n38899), .B1(n5019), .B2(n35677), .ZN(
        n7186) );
  OAI22_X1 U1471 ( .A1(n37975), .A2(n38850), .B1(n4948), .B2(n35857), .ZN(
        n7243) );
  OAI22_X1 U1472 ( .A1(n37976), .A2(n38857), .B1(n4948), .B2(n35866), .ZN(
        n7244) );
  OAI22_X1 U1473 ( .A1(n37976), .A2(n38864), .B1(n4948), .B2(n35875), .ZN(
        n7245) );
  OAI22_X1 U1474 ( .A1(n37976), .A2(n38871), .B1(n37970), .B2(n35884), .ZN(
        n7246) );
  OAI22_X1 U1475 ( .A1(n37976), .A2(n38878), .B1(n37970), .B2(n35893), .ZN(
        n7247) );
  OAI22_X1 U1476 ( .A1(n37976), .A2(n38885), .B1(n37970), .B2(n35902), .ZN(
        n7248) );
  OAI22_X1 U1477 ( .A1(n37977), .A2(n38892), .B1(n37970), .B2(n35911), .ZN(
        n7249) );
  OAI22_X1 U1478 ( .A1(n37977), .A2(n38899), .B1(n4948), .B2(n35920), .ZN(
        n7250) );
  OAI22_X1 U1479 ( .A1(n37987), .A2(n38850), .B1(n4913), .B2(n35346), .ZN(
        n7275) );
  OAI22_X1 U1480 ( .A1(n37988), .A2(n38857), .B1(n4913), .B2(n35355), .ZN(
        n7276) );
  OAI22_X1 U1481 ( .A1(n37988), .A2(n38864), .B1(n4913), .B2(n35364), .ZN(
        n7277) );
  OAI22_X1 U1482 ( .A1(n37988), .A2(n38871), .B1(n37982), .B2(n35373), .ZN(
        n7278) );
  OAI22_X1 U1483 ( .A1(n37988), .A2(n38878), .B1(n37982), .B2(n35382), .ZN(
        n7279) );
  OAI22_X1 U1484 ( .A1(n37988), .A2(n38885), .B1(n37982), .B2(n35391), .ZN(
        n7280) );
  OAI22_X1 U1485 ( .A1(n37989), .A2(n38892), .B1(n37982), .B2(n35400), .ZN(
        n7281) );
  OAI22_X1 U1486 ( .A1(n37989), .A2(n38899), .B1(n4913), .B2(n35409), .ZN(
        n7282) );
  OAI22_X1 U1487 ( .A1(n38008), .A2(n38850), .B1(n4843), .B2(n36367), .ZN(
        n7339) );
  OAI22_X1 U1488 ( .A1(n38009), .A2(n38857), .B1(n4843), .B2(n36376), .ZN(
        n7340) );
  OAI22_X1 U1489 ( .A1(n38009), .A2(n38864), .B1(n4843), .B2(n36385), .ZN(
        n7341) );
  OAI22_X1 U1490 ( .A1(n38009), .A2(n38871), .B1(n38003), .B2(n36394), .ZN(
        n7342) );
  OAI22_X1 U1491 ( .A1(n38009), .A2(n38878), .B1(n38003), .B2(n36403), .ZN(
        n7343) );
  OAI22_X1 U1492 ( .A1(n38009), .A2(n38885), .B1(n38003), .B2(n36412), .ZN(
        n7344) );
  OAI22_X1 U1493 ( .A1(n38010), .A2(n38892), .B1(n38003), .B2(n36421), .ZN(
        n7345) );
  OAI22_X1 U1494 ( .A1(n38010), .A2(n38899), .B1(n4843), .B2(n36430), .ZN(
        n7346) );
  OAI22_X1 U1495 ( .A1(n38029), .A2(n38850), .B1(n4773), .B2(n35856), .ZN(
        n7403) );
  OAI22_X1 U1496 ( .A1(n38030), .A2(n38857), .B1(n4773), .B2(n35865), .ZN(
        n7404) );
  OAI22_X1 U1497 ( .A1(n38030), .A2(n38864), .B1(n4773), .B2(n35874), .ZN(
        n7405) );
  OAI22_X1 U1498 ( .A1(n38030), .A2(n38871), .B1(n38024), .B2(n35883), .ZN(
        n7406) );
  OAI22_X1 U1499 ( .A1(n38030), .A2(n38878), .B1(n38024), .B2(n35892), .ZN(
        n7407) );
  OAI22_X1 U1500 ( .A1(n38030), .A2(n38885), .B1(n38024), .B2(n35901), .ZN(
        n7408) );
  OAI22_X1 U1501 ( .A1(n38031), .A2(n38892), .B1(n38024), .B2(n35910), .ZN(
        n7409) );
  OAI22_X1 U1502 ( .A1(n38031), .A2(n38899), .B1(n4773), .B2(n35919), .ZN(
        n7410) );
  OAI22_X1 U1503 ( .A1(n38041), .A2(n38850), .B1(n4738), .B2(n35349), .ZN(
        n7435) );
  OAI22_X1 U1504 ( .A1(n38042), .A2(n38857), .B1(n4738), .B2(n35358), .ZN(
        n7436) );
  OAI22_X1 U1505 ( .A1(n38042), .A2(n38864), .B1(n4738), .B2(n35367), .ZN(
        n7437) );
  OAI22_X1 U1506 ( .A1(n38042), .A2(n38871), .B1(n38036), .B2(n35376), .ZN(
        n7438) );
  OAI22_X1 U1507 ( .A1(n38042), .A2(n38878), .B1(n38036), .B2(n35385), .ZN(
        n7439) );
  OAI22_X1 U1508 ( .A1(n38042), .A2(n38885), .B1(n38036), .B2(n35394), .ZN(
        n7440) );
  OAI22_X1 U1509 ( .A1(n38043), .A2(n38892), .B1(n38036), .B2(n35403), .ZN(
        n7441) );
  OAI22_X1 U1510 ( .A1(n38043), .A2(n38899), .B1(n4738), .B2(n35412), .ZN(
        n7442) );
  OAI22_X1 U1511 ( .A1(n38062), .A2(n38850), .B1(n4668), .B2(n36374), .ZN(
        n7499) );
  OAI22_X1 U1512 ( .A1(n38063), .A2(n38857), .B1(n4668), .B2(n36383), .ZN(
        n7500) );
  OAI22_X1 U1513 ( .A1(n38063), .A2(n38864), .B1(n4668), .B2(n36392), .ZN(
        n7501) );
  OAI22_X1 U1514 ( .A1(n38063), .A2(n38871), .B1(n38057), .B2(n36401), .ZN(
        n7502) );
  OAI22_X1 U1515 ( .A1(n38063), .A2(n38878), .B1(n38057), .B2(n36410), .ZN(
        n7503) );
  OAI22_X1 U1516 ( .A1(n38063), .A2(n38885), .B1(n38057), .B2(n36419), .ZN(
        n7504) );
  OAI22_X1 U1517 ( .A1(n38064), .A2(n38892), .B1(n38057), .B2(n36428), .ZN(
        n7505) );
  OAI22_X1 U1518 ( .A1(n38064), .A2(n38899), .B1(n4668), .B2(n36437), .ZN(
        n7506) );
  OAI22_X1 U1519 ( .A1(n38083), .A2(n38849), .B1(n4598), .B2(n35859), .ZN(
        n7563) );
  OAI22_X1 U1520 ( .A1(n38084), .A2(n38856), .B1(n4598), .B2(n35868), .ZN(
        n7564) );
  OAI22_X1 U1521 ( .A1(n38084), .A2(n38863), .B1(n4598), .B2(n35877), .ZN(
        n7565) );
  OAI22_X1 U1522 ( .A1(n38084), .A2(n38870), .B1(n38078), .B2(n35886), .ZN(
        n7566) );
  OAI22_X1 U1523 ( .A1(n38084), .A2(n38877), .B1(n38078), .B2(n35895), .ZN(
        n7567) );
  OAI22_X1 U1524 ( .A1(n38084), .A2(n38884), .B1(n38078), .B2(n35904), .ZN(
        n7568) );
  OAI22_X1 U1525 ( .A1(n38085), .A2(n38891), .B1(n38078), .B2(n35913), .ZN(
        n7569) );
  OAI22_X1 U1526 ( .A1(n38085), .A2(n38898), .B1(n4598), .B2(n35922), .ZN(
        n7570) );
  OAI22_X1 U1527 ( .A1(n38095), .A2(n38849), .B1(n4563), .B2(n35348), .ZN(
        n7595) );
  OAI22_X1 U1528 ( .A1(n38096), .A2(n38856), .B1(n4563), .B2(n35357), .ZN(
        n7596) );
  OAI22_X1 U1529 ( .A1(n38096), .A2(n38863), .B1(n4563), .B2(n35366), .ZN(
        n7597) );
  OAI22_X1 U1530 ( .A1(n38096), .A2(n38870), .B1(n38090), .B2(n35375), .ZN(
        n7598) );
  OAI22_X1 U1531 ( .A1(n38096), .A2(n38877), .B1(n38090), .B2(n35384), .ZN(
        n7599) );
  OAI22_X1 U1532 ( .A1(n38096), .A2(n38884), .B1(n38090), .B2(n35393), .ZN(
        n7600) );
  OAI22_X1 U1533 ( .A1(n38097), .A2(n38891), .B1(n38090), .B2(n35402), .ZN(
        n7601) );
  OAI22_X1 U1534 ( .A1(n38097), .A2(n38898), .B1(n4563), .B2(n35411), .ZN(
        n7602) );
  OAI22_X1 U1535 ( .A1(n38116), .A2(n38849), .B1(n4493), .B2(n36190), .ZN(
        n7659) );
  OAI22_X1 U1536 ( .A1(n38117), .A2(n38856), .B1(n4493), .B2(n36191), .ZN(
        n7660) );
  OAI22_X1 U1537 ( .A1(n38117), .A2(n38863), .B1(n4493), .B2(n36192), .ZN(
        n7661) );
  OAI22_X1 U1538 ( .A1(n38117), .A2(n38870), .B1(n38111), .B2(n36193), .ZN(
        n7662) );
  OAI22_X1 U1539 ( .A1(n38117), .A2(n38877), .B1(n38111), .B2(n36194), .ZN(
        n7663) );
  OAI22_X1 U1540 ( .A1(n38117), .A2(n38884), .B1(n38111), .B2(n36195), .ZN(
        n7664) );
  OAI22_X1 U1541 ( .A1(n38118), .A2(n38891), .B1(n38111), .B2(n36196), .ZN(
        n7665) );
  OAI22_X1 U1542 ( .A1(n38118), .A2(n38898), .B1(n4493), .B2(n36197), .ZN(
        n7666) );
  OAI22_X1 U1543 ( .A1(n38137), .A2(n38849), .B1(n4423), .B2(n35678), .ZN(
        n7723) );
  OAI22_X1 U1544 ( .A1(n38138), .A2(n38856), .B1(n4423), .B2(n35679), .ZN(
        n7724) );
  OAI22_X1 U1545 ( .A1(n38138), .A2(n38863), .B1(n4423), .B2(n35680), .ZN(
        n7725) );
  OAI22_X1 U1546 ( .A1(n38138), .A2(n38870), .B1(n38132), .B2(n35681), .ZN(
        n7726) );
  OAI22_X1 U1547 ( .A1(n38138), .A2(n38877), .B1(n38132), .B2(n35682), .ZN(
        n7727) );
  OAI22_X1 U1548 ( .A1(n38138), .A2(n38884), .B1(n38132), .B2(n35683), .ZN(
        n7728) );
  OAI22_X1 U1549 ( .A1(n38139), .A2(n38891), .B1(n38132), .B2(n35684), .ZN(
        n7729) );
  OAI22_X1 U1550 ( .A1(n38139), .A2(n38898), .B1(n4423), .B2(n35685), .ZN(
        n7730) );
  OAI22_X1 U1551 ( .A1(n38149), .A2(n38849), .B1(n4388), .B2(n36369), .ZN(
        n7755) );
  OAI22_X1 U1552 ( .A1(n38150), .A2(n38856), .B1(n4388), .B2(n36378), .ZN(
        n7756) );
  OAI22_X1 U1553 ( .A1(n38150), .A2(n38863), .B1(n4388), .B2(n36387), .ZN(
        n7757) );
  OAI22_X1 U1554 ( .A1(n38150), .A2(n38870), .B1(n38144), .B2(n36396), .ZN(
        n7758) );
  OAI22_X1 U1555 ( .A1(n38150), .A2(n38877), .B1(n38144), .B2(n36405), .ZN(
        n7759) );
  OAI22_X1 U1556 ( .A1(n38150), .A2(n38884), .B1(n38144), .B2(n36414), .ZN(
        n7760) );
  OAI22_X1 U1557 ( .A1(n38151), .A2(n38891), .B1(n38144), .B2(n36423), .ZN(
        n7761) );
  OAI22_X1 U1558 ( .A1(n38151), .A2(n38898), .B1(n4388), .B2(n36432), .ZN(
        n7762) );
  OAI22_X1 U1559 ( .A1(n38170), .A2(n38849), .B1(n4318), .B2(n35858), .ZN(
        n7819) );
  OAI22_X1 U1560 ( .A1(n38171), .A2(n38856), .B1(n4318), .B2(n35867), .ZN(
        n7820) );
  OAI22_X1 U1561 ( .A1(n38171), .A2(n38863), .B1(n4318), .B2(n35876), .ZN(
        n7821) );
  OAI22_X1 U1562 ( .A1(n38171), .A2(n38870), .B1(n38165), .B2(n35885), .ZN(
        n7822) );
  OAI22_X1 U1563 ( .A1(n38171), .A2(n38877), .B1(n38165), .B2(n35894), .ZN(
        n7823) );
  OAI22_X1 U1564 ( .A1(n38171), .A2(n38884), .B1(n38165), .B2(n35903), .ZN(
        n7824) );
  OAI22_X1 U1565 ( .A1(n38172), .A2(n38891), .B1(n38165), .B2(n35912), .ZN(
        n7825) );
  OAI22_X1 U1566 ( .A1(n38172), .A2(n38898), .B1(n4318), .B2(n35921), .ZN(
        n7826) );
  OAI22_X1 U1567 ( .A1(n38182), .A2(n38849), .B1(n4283), .B2(n35343), .ZN(
        n7851) );
  OAI22_X1 U1568 ( .A1(n38183), .A2(n38856), .B1(n4283), .B2(n35352), .ZN(
        n7852) );
  OAI22_X1 U1569 ( .A1(n38183), .A2(n38863), .B1(n4283), .B2(n35361), .ZN(
        n7853) );
  OAI22_X1 U1570 ( .A1(n38183), .A2(n38870), .B1(n38177), .B2(n35370), .ZN(
        n7854) );
  OAI22_X1 U1571 ( .A1(n38183), .A2(n38877), .B1(n38177), .B2(n35379), .ZN(
        n7855) );
  OAI22_X1 U1572 ( .A1(n38183), .A2(n38884), .B1(n38177), .B2(n35388), .ZN(
        n7856) );
  OAI22_X1 U1573 ( .A1(n38184), .A2(n38891), .B1(n38177), .B2(n35397), .ZN(
        n7857) );
  OAI22_X1 U1574 ( .A1(n38184), .A2(n38898), .B1(n4283), .B2(n35406), .ZN(
        n7858) );
  OAI22_X1 U1575 ( .A1(n38203), .A2(n38848), .B1(n4213), .B2(n36368), .ZN(
        n7915) );
  OAI22_X1 U1576 ( .A1(n38204), .A2(n38855), .B1(n4213), .B2(n36377), .ZN(
        n7916) );
  OAI22_X1 U1577 ( .A1(n38204), .A2(n38862), .B1(n4213), .B2(n36386), .ZN(
        n7917) );
  OAI22_X1 U1578 ( .A1(n38204), .A2(n38869), .B1(n38198), .B2(n36395), .ZN(
        n7918) );
  OAI22_X1 U1579 ( .A1(n38204), .A2(n38876), .B1(n38198), .B2(n36404), .ZN(
        n7919) );
  OAI22_X1 U1580 ( .A1(n38204), .A2(n38883), .B1(n38198), .B2(n36413), .ZN(
        n7920) );
  OAI22_X1 U1581 ( .A1(n38205), .A2(n38890), .B1(n38198), .B2(n36422), .ZN(
        n7921) );
  OAI22_X1 U1582 ( .A1(n38205), .A2(n38897), .B1(n4213), .B2(n36431), .ZN(
        n7922) );
  OAI22_X1 U1583 ( .A1(n38224), .A2(n38848), .B1(n4140), .B2(n35861), .ZN(
        n7979) );
  OAI22_X1 U1584 ( .A1(n38225), .A2(n38855), .B1(n4140), .B2(n35870), .ZN(
        n7980) );
  OAI22_X1 U1585 ( .A1(n38225), .A2(n38862), .B1(n4140), .B2(n35879), .ZN(
        n7981) );
  OAI22_X1 U1586 ( .A1(n38225), .A2(n38869), .B1(n38219), .B2(n35888), .ZN(
        n7982) );
  OAI22_X1 U1587 ( .A1(n38225), .A2(n38876), .B1(n38219), .B2(n35897), .ZN(
        n7983) );
  OAI22_X1 U1588 ( .A1(n38225), .A2(n38883), .B1(n38219), .B2(n35906), .ZN(
        n7984) );
  OAI22_X1 U1589 ( .A1(n38226), .A2(n38890), .B1(n38219), .B2(n35915), .ZN(
        n7985) );
  OAI22_X1 U1590 ( .A1(n38226), .A2(n38897), .B1(n4140), .B2(n35924), .ZN(
        n7986) );
  OAI22_X1 U1591 ( .A1(n38236), .A2(n38848), .B1(n4076), .B2(n35350), .ZN(
        n8011) );
  OAI22_X1 U1592 ( .A1(n38237), .A2(n38855), .B1(n4076), .B2(n35359), .ZN(
        n8012) );
  OAI22_X1 U1593 ( .A1(n38237), .A2(n38862), .B1(n4076), .B2(n35368), .ZN(
        n8013) );
  OAI22_X1 U1594 ( .A1(n38237), .A2(n38869), .B1(n38231), .B2(n35377), .ZN(
        n8014) );
  OAI22_X1 U1595 ( .A1(n38237), .A2(n38876), .B1(n38231), .B2(n35386), .ZN(
        n8015) );
  OAI22_X1 U1596 ( .A1(n38237), .A2(n38883), .B1(n38231), .B2(n35395), .ZN(
        n8016) );
  OAI22_X1 U1597 ( .A1(n38238), .A2(n38890), .B1(n38231), .B2(n35404), .ZN(
        n8017) );
  OAI22_X1 U1598 ( .A1(n38238), .A2(n38897), .B1(n4076), .B2(n35413), .ZN(
        n8018) );
  OAI22_X1 U1599 ( .A1(n38257), .A2(n38848), .B1(n4006), .B2(n36371), .ZN(
        n8075) );
  OAI22_X1 U1600 ( .A1(n38258), .A2(n38855), .B1(n4006), .B2(n36380), .ZN(
        n8076) );
  OAI22_X1 U1601 ( .A1(n38258), .A2(n38862), .B1(n4006), .B2(n36389), .ZN(
        n8077) );
  OAI22_X1 U1602 ( .A1(n38258), .A2(n38869), .B1(n38252), .B2(n36398), .ZN(
        n8078) );
  OAI22_X1 U1603 ( .A1(n38258), .A2(n38876), .B1(n38252), .B2(n36407), .ZN(
        n8079) );
  OAI22_X1 U1604 ( .A1(n38258), .A2(n38883), .B1(n38252), .B2(n36416), .ZN(
        n8080) );
  OAI22_X1 U1605 ( .A1(n38259), .A2(n38890), .B1(n38252), .B2(n36425), .ZN(
        n8081) );
  OAI22_X1 U1606 ( .A1(n38259), .A2(n38897), .B1(n4006), .B2(n36434), .ZN(
        n8082) );
  OAI22_X1 U1607 ( .A1(n38278), .A2(n38848), .B1(n3936), .B2(n35860), .ZN(
        n8139) );
  OAI22_X1 U1608 ( .A1(n38279), .A2(n38855), .B1(n3936), .B2(n35869), .ZN(
        n8140) );
  OAI22_X1 U1609 ( .A1(n38279), .A2(n38862), .B1(n3936), .B2(n35878), .ZN(
        n8141) );
  OAI22_X1 U1610 ( .A1(n38279), .A2(n38869), .B1(n38273), .B2(n35887), .ZN(
        n8142) );
  OAI22_X1 U1611 ( .A1(n38279), .A2(n38876), .B1(n38273), .B2(n35896), .ZN(
        n8143) );
  OAI22_X1 U1612 ( .A1(n38279), .A2(n38883), .B1(n38273), .B2(n35905), .ZN(
        n8144) );
  OAI22_X1 U1613 ( .A1(n38280), .A2(n38890), .B1(n38273), .B2(n35914), .ZN(
        n8145) );
  OAI22_X1 U1614 ( .A1(n38280), .A2(n38897), .B1(n3936), .B2(n35923), .ZN(
        n8146) );
  OAI22_X1 U1615 ( .A1(n38290), .A2(n38848), .B1(n3901), .B2(n35166), .ZN(
        n8171) );
  OAI22_X1 U1616 ( .A1(n38291), .A2(n38855), .B1(n3901), .B2(n35167), .ZN(
        n8172) );
  OAI22_X1 U1617 ( .A1(n38291), .A2(n38862), .B1(n3901), .B2(n35168), .ZN(
        n8173) );
  OAI22_X1 U1618 ( .A1(n38291), .A2(n38869), .B1(n38285), .B2(n35169), .ZN(
        n8174) );
  OAI22_X1 U1619 ( .A1(n38291), .A2(n38876), .B1(n38285), .B2(n35170), .ZN(
        n8175) );
  OAI22_X1 U1620 ( .A1(n38291), .A2(n38883), .B1(n38285), .B2(n35171), .ZN(
        n8176) );
  OAI22_X1 U1621 ( .A1(n38292), .A2(n38890), .B1(n38285), .B2(n35172), .ZN(
        n8177) );
  OAI22_X1 U1622 ( .A1(n38292), .A2(n38897), .B1(n3901), .B2(n35173), .ZN(
        n8178) );
  OAI22_X1 U1623 ( .A1(n38311), .A2(n38848), .B1(n3831), .B2(n36198), .ZN(
        n8235) );
  OAI22_X1 U1624 ( .A1(n38312), .A2(n38855), .B1(n3831), .B2(n36199), .ZN(
        n8236) );
  OAI22_X1 U1625 ( .A1(n38312), .A2(n38862), .B1(n3831), .B2(n36200), .ZN(
        n8237) );
  OAI22_X1 U1626 ( .A1(n38312), .A2(n38869), .B1(n38306), .B2(n36201), .ZN(
        n8238) );
  OAI22_X1 U1627 ( .A1(n38312), .A2(n38876), .B1(n38306), .B2(n36202), .ZN(
        n8239) );
  OAI22_X1 U1628 ( .A1(n38312), .A2(n38883), .B1(n38306), .B2(n36203), .ZN(
        n8240) );
  OAI22_X1 U1629 ( .A1(n38313), .A2(n38890), .B1(n38306), .B2(n36204), .ZN(
        n8241) );
  OAI22_X1 U1630 ( .A1(n38313), .A2(n38897), .B1(n3831), .B2(n36205), .ZN(
        n8242) );
  OAI22_X1 U1631 ( .A1(n38323), .A2(n38848), .B1(n3796), .B2(n35345), .ZN(
        n8267) );
  OAI22_X1 U1632 ( .A1(n38324), .A2(n38855), .B1(n3796), .B2(n35354), .ZN(
        n8268) );
  OAI22_X1 U1633 ( .A1(n38324), .A2(n38862), .B1(n3796), .B2(n35363), .ZN(
        n8269) );
  OAI22_X1 U1634 ( .A1(n38324), .A2(n38869), .B1(n38318), .B2(n35372), .ZN(
        n8270) );
  OAI22_X1 U1635 ( .A1(n38324), .A2(n38876), .B1(n38318), .B2(n35381), .ZN(
        n8271) );
  OAI22_X1 U1636 ( .A1(n38324), .A2(n38883), .B1(n38318), .B2(n35390), .ZN(
        n8272) );
  OAI22_X1 U1637 ( .A1(n38325), .A2(n38890), .B1(n38318), .B2(n35399), .ZN(
        n8273) );
  OAI22_X1 U1638 ( .A1(n38325), .A2(n38897), .B1(n3796), .B2(n35408), .ZN(
        n8274) );
  OAI22_X1 U1639 ( .A1(n38344), .A2(n38847), .B1(n3726), .B2(n36370), .ZN(
        n8331) );
  OAI22_X1 U1640 ( .A1(n38345), .A2(n38854), .B1(n3726), .B2(n36379), .ZN(
        n8332) );
  OAI22_X1 U1641 ( .A1(n38345), .A2(n38861), .B1(n3726), .B2(n36388), .ZN(
        n8333) );
  OAI22_X1 U1642 ( .A1(n38345), .A2(n38868), .B1(n38339), .B2(n36397), .ZN(
        n8334) );
  OAI22_X1 U1643 ( .A1(n38345), .A2(n38875), .B1(n38339), .B2(n36406), .ZN(
        n8335) );
  OAI22_X1 U1644 ( .A1(n38345), .A2(n38882), .B1(n38339), .B2(n36415), .ZN(
        n8336) );
  OAI22_X1 U1645 ( .A1(n38346), .A2(n38889), .B1(n38339), .B2(n36424), .ZN(
        n8337) );
  OAI22_X1 U1646 ( .A1(n38346), .A2(n38896), .B1(n3726), .B2(n36433), .ZN(
        n8338) );
  OAI22_X1 U1647 ( .A1(n38365), .A2(n38847), .B1(n3656), .B2(n35855), .ZN(
        n8395) );
  OAI22_X1 U1648 ( .A1(n38366), .A2(n38854), .B1(n3656), .B2(n35864), .ZN(
        n8396) );
  OAI22_X1 U1649 ( .A1(n38366), .A2(n38861), .B1(n3656), .B2(n35873), .ZN(
        n8397) );
  OAI22_X1 U1650 ( .A1(n38366), .A2(n38868), .B1(n38360), .B2(n35882), .ZN(
        n8398) );
  OAI22_X1 U1651 ( .A1(n38366), .A2(n38875), .B1(n38360), .B2(n35891), .ZN(
        n8399) );
  OAI22_X1 U1652 ( .A1(n38366), .A2(n38882), .B1(n38360), .B2(n35900), .ZN(
        n8400) );
  OAI22_X1 U1653 ( .A1(n38367), .A2(n38889), .B1(n38360), .B2(n35909), .ZN(
        n8401) );
  OAI22_X1 U1654 ( .A1(n38367), .A2(n38896), .B1(n3656), .B2(n35918), .ZN(
        n8402) );
  OAI22_X1 U1655 ( .A1(n38377), .A2(n38847), .B1(n3621), .B2(n35344), .ZN(
        n8427) );
  OAI22_X1 U1656 ( .A1(n38378), .A2(n38854), .B1(n3621), .B2(n35353), .ZN(
        n8428) );
  OAI22_X1 U1657 ( .A1(n38378), .A2(n38861), .B1(n3621), .B2(n35362), .ZN(
        n8429) );
  OAI22_X1 U1658 ( .A1(n38378), .A2(n38868), .B1(n38372), .B2(n35371), .ZN(
        n8430) );
  OAI22_X1 U1659 ( .A1(n38378), .A2(n38875), .B1(n38372), .B2(n35380), .ZN(
        n8431) );
  OAI22_X1 U1660 ( .A1(n38378), .A2(n38882), .B1(n38372), .B2(n35389), .ZN(
        n8432) );
  OAI22_X1 U1661 ( .A1(n38379), .A2(n38889), .B1(n38372), .B2(n35398), .ZN(
        n8433) );
  OAI22_X1 U1662 ( .A1(n38379), .A2(n38896), .B1(n3621), .B2(n35407), .ZN(
        n8434) );
  OAI22_X1 U1663 ( .A1(n38398), .A2(n38847), .B1(n3551), .B2(n36373), .ZN(
        n8491) );
  OAI22_X1 U1664 ( .A1(n38399), .A2(n38854), .B1(n3551), .B2(n36382), .ZN(
        n8492) );
  OAI22_X1 U1665 ( .A1(n38399), .A2(n38861), .B1(n3551), .B2(n36391), .ZN(
        n8493) );
  OAI22_X1 U1666 ( .A1(n38399), .A2(n38868), .B1(n38393), .B2(n36400), .ZN(
        n8494) );
  OAI22_X1 U1667 ( .A1(n38399), .A2(n38875), .B1(n38393), .B2(n36409), .ZN(
        n8495) );
  OAI22_X1 U1668 ( .A1(n38399), .A2(n38882), .B1(n38393), .B2(n36418), .ZN(
        n8496) );
  OAI22_X1 U1669 ( .A1(n38400), .A2(n38889), .B1(n38393), .B2(n36427), .ZN(
        n8497) );
  OAI22_X1 U1670 ( .A1(n38400), .A2(n38896), .B1(n3551), .B2(n36436), .ZN(
        n8498) );
  OAI22_X1 U1671 ( .A1(n38419), .A2(n38847), .B1(n3481), .B2(n35862), .ZN(
        n8555) );
  OAI22_X1 U1672 ( .A1(n38420), .A2(n38854), .B1(n3481), .B2(n35871), .ZN(
        n8556) );
  OAI22_X1 U1673 ( .A1(n38420), .A2(n38861), .B1(n3481), .B2(n35880), .ZN(
        n8557) );
  OAI22_X1 U1674 ( .A1(n38420), .A2(n38868), .B1(n38414), .B2(n35889), .ZN(
        n8558) );
  OAI22_X1 U1675 ( .A1(n38420), .A2(n38875), .B1(n38414), .B2(n35898), .ZN(
        n8559) );
  OAI22_X1 U1676 ( .A1(n38420), .A2(n38882), .B1(n38414), .B2(n35907), .ZN(
        n8560) );
  OAI22_X1 U1677 ( .A1(n38421), .A2(n38889), .B1(n38414), .B2(n35916), .ZN(
        n8561) );
  OAI22_X1 U1678 ( .A1(n38421), .A2(n38896), .B1(n3481), .B2(n35925), .ZN(
        n8562) );
  OAI22_X1 U1679 ( .A1(n38431), .A2(n38847), .B1(n3446), .B2(n35347), .ZN(
        n8587) );
  OAI22_X1 U1680 ( .A1(n38432), .A2(n38854), .B1(n3446), .B2(n35356), .ZN(
        n8588) );
  OAI22_X1 U1681 ( .A1(n38432), .A2(n38861), .B1(n3446), .B2(n35365), .ZN(
        n8589) );
  OAI22_X1 U1682 ( .A1(n38432), .A2(n38868), .B1(n38426), .B2(n35374), .ZN(
        n8590) );
  OAI22_X1 U1683 ( .A1(n38432), .A2(n38875), .B1(n38426), .B2(n35383), .ZN(
        n8591) );
  OAI22_X1 U1684 ( .A1(n38432), .A2(n38882), .B1(n38426), .B2(n35392), .ZN(
        n8592) );
  OAI22_X1 U1685 ( .A1(n38433), .A2(n38889), .B1(n38426), .B2(n35401), .ZN(
        n8593) );
  OAI22_X1 U1686 ( .A1(n38433), .A2(n38896), .B1(n3446), .B2(n35410), .ZN(
        n8594) );
  OAI22_X1 U1687 ( .A1(n38452), .A2(n38847), .B1(n3376), .B2(n36372), .ZN(
        n8651) );
  OAI22_X1 U1688 ( .A1(n38453), .A2(n38854), .B1(n3376), .B2(n36381), .ZN(
        n8652) );
  OAI22_X1 U1689 ( .A1(n38453), .A2(n38861), .B1(n3376), .B2(n36390), .ZN(
        n8653) );
  OAI22_X1 U1690 ( .A1(n38453), .A2(n38868), .B1(n38447), .B2(n36399), .ZN(
        n8654) );
  OAI22_X1 U1691 ( .A1(n38453), .A2(n38875), .B1(n38447), .B2(n36408), .ZN(
        n8655) );
  OAI22_X1 U1692 ( .A1(n38453), .A2(n38882), .B1(n38447), .B2(n36417), .ZN(
        n8656) );
  OAI22_X1 U1693 ( .A1(n38454), .A2(n38889), .B1(n38447), .B2(n36426), .ZN(
        n8657) );
  OAI22_X1 U1694 ( .A1(n38454), .A2(n38896), .B1(n3376), .B2(n36435), .ZN(
        n8658) );
  OAI22_X1 U1695 ( .A1(n38473), .A2(n38846), .B1(n3306), .B2(n35686), .ZN(
        n8715) );
  OAI22_X1 U1696 ( .A1(n38474), .A2(n38853), .B1(n3306), .B2(n35687), .ZN(
        n8716) );
  OAI22_X1 U1697 ( .A1(n38474), .A2(n38860), .B1(n3306), .B2(n35688), .ZN(
        n8717) );
  OAI22_X1 U1698 ( .A1(n38474), .A2(n38867), .B1(n38468), .B2(n35689), .ZN(
        n8718) );
  OAI22_X1 U1699 ( .A1(n38474), .A2(n38874), .B1(n38468), .B2(n35690), .ZN(
        n8719) );
  OAI22_X1 U1700 ( .A1(n38474), .A2(n38881), .B1(n38468), .B2(n35691), .ZN(
        n8720) );
  OAI22_X1 U1701 ( .A1(n38475), .A2(n38888), .B1(n38468), .B2(n35692), .ZN(
        n8721) );
  OAI22_X1 U1702 ( .A1(n38475), .A2(n38895), .B1(n3306), .B2(n35693), .ZN(
        n8722) );
  OAI22_X1 U1703 ( .A1(n38491), .A2(n38846), .B1(n3270), .B2(n35174), .ZN(
        n8747) );
  OAI22_X1 U1704 ( .A1(n38492), .A2(n38853), .B1(n3270), .B2(n35175), .ZN(
        n8748) );
  OAI22_X1 U1705 ( .A1(n38492), .A2(n38860), .B1(n3270), .B2(n35176), .ZN(
        n8749) );
  OAI22_X1 U1706 ( .A1(n38492), .A2(n38867), .B1(n38486), .B2(n35177), .ZN(
        n8750) );
  OAI22_X1 U1707 ( .A1(n38492), .A2(n38874), .B1(n38486), .B2(n35178), .ZN(
        n8751) );
  OAI22_X1 U1708 ( .A1(n38492), .A2(n38881), .B1(n38486), .B2(n35179), .ZN(
        n8752) );
  OAI22_X1 U1709 ( .A1(n38493), .A2(n38888), .B1(n38486), .B2(n35180), .ZN(
        n8753) );
  OAI22_X1 U1710 ( .A1(n38493), .A2(n38895), .B1(n3270), .B2(n35181), .ZN(
        n8754) );
  OAI22_X1 U1711 ( .A1(n38515), .A2(n38846), .B1(n3200), .B2(n35182), .ZN(
        n8811) );
  OAI22_X1 U1712 ( .A1(n38516), .A2(n38853), .B1(n38510), .B2(n35183), .ZN(
        n8812) );
  OAI22_X1 U1713 ( .A1(n38516), .A2(n38860), .B1(n38510), .B2(n35184), .ZN(
        n8813) );
  OAI22_X1 U1714 ( .A1(n38516), .A2(n38867), .B1(n38510), .B2(n35185), .ZN(
        n8814) );
  OAI22_X1 U1715 ( .A1(n38516), .A2(n38874), .B1(n38510), .B2(n35186), .ZN(
        n8815) );
  OAI22_X1 U1716 ( .A1(n38516), .A2(n38881), .B1(n38510), .B2(n35187), .ZN(
        n8816) );
  OAI22_X1 U1717 ( .A1(n38517), .A2(n38888), .B1(n38510), .B2(n35188), .ZN(
        n8817) );
  OAI22_X1 U1718 ( .A1(n38517), .A2(n38895), .B1(n3200), .B2(n35189), .ZN(
        n8818) );
  OAI22_X1 U1719 ( .A1(n38527), .A2(n38846), .B1(n3165), .B2(n36206), .ZN(
        n8843) );
  OAI22_X1 U1720 ( .A1(n38528), .A2(n38853), .B1(n38522), .B2(n36207), .ZN(
        n8844) );
  OAI22_X1 U1721 ( .A1(n38528), .A2(n38860), .B1(n38522), .B2(n36208), .ZN(
        n8845) );
  OAI22_X1 U1722 ( .A1(n38528), .A2(n38867), .B1(n38522), .B2(n36209), .ZN(
        n8846) );
  OAI22_X1 U1723 ( .A1(n38528), .A2(n38874), .B1(n38522), .B2(n36210), .ZN(
        n8847) );
  OAI22_X1 U1724 ( .A1(n38528), .A2(n38881), .B1(n38522), .B2(n36211), .ZN(
        n8848) );
  OAI22_X1 U1725 ( .A1(n38529), .A2(n38888), .B1(n38522), .B2(n36212), .ZN(
        n8849) );
  OAI22_X1 U1726 ( .A1(n38529), .A2(n38895), .B1(n3165), .B2(n36213), .ZN(
        n8850) );
  OAI22_X1 U1727 ( .A1(n38539), .A2(n38846), .B1(n3130), .B2(n35694), .ZN(
        n8875) );
  OAI22_X1 U1728 ( .A1(n38540), .A2(n38853), .B1(n38534), .B2(n35695), .ZN(
        n8876) );
  OAI22_X1 U1729 ( .A1(n38540), .A2(n38860), .B1(n38534), .B2(n35696), .ZN(
        n8877) );
  OAI22_X1 U1730 ( .A1(n38540), .A2(n38867), .B1(n38534), .B2(n35697), .ZN(
        n8878) );
  OAI22_X1 U1731 ( .A1(n38540), .A2(n38874), .B1(n38534), .B2(n35698), .ZN(
        n8879) );
  OAI22_X1 U1732 ( .A1(n38540), .A2(n38881), .B1(n38534), .B2(n35699), .ZN(
        n8880) );
  OAI22_X1 U1733 ( .A1(n38541), .A2(n38888), .B1(n38534), .B2(n35700), .ZN(
        n8881) );
  OAI22_X1 U1734 ( .A1(n38541), .A2(n38895), .B1(n3130), .B2(n35701), .ZN(
        n8882) );
  OAI22_X1 U1735 ( .A1(n38575), .A2(n38846), .B1(n3025), .B2(n35510), .ZN(
        n8971) );
  OAI22_X1 U1736 ( .A1(n38576), .A2(n38853), .B1(n38570), .B2(n35511), .ZN(
        n8972) );
  OAI22_X1 U1737 ( .A1(n38576), .A2(n38860), .B1(n38570), .B2(n35512), .ZN(
        n8973) );
  OAI22_X1 U1738 ( .A1(n38576), .A2(n38867), .B1(n38570), .B2(n35513), .ZN(
        n8974) );
  OAI22_X1 U1739 ( .A1(n38576), .A2(n38874), .B1(n38570), .B2(n35514), .ZN(
        n8975) );
  OAI22_X1 U1740 ( .A1(n38576), .A2(n38881), .B1(n38570), .B2(n35515), .ZN(
        n8976) );
  OAI22_X1 U1741 ( .A1(n38577), .A2(n38888), .B1(n38570), .B2(n35516), .ZN(
        n8977) );
  OAI22_X1 U1742 ( .A1(n38577), .A2(n38895), .B1(n3025), .B2(n35517), .ZN(
        n8978) );
  OAI22_X1 U1743 ( .A1(n38587), .A2(n38846), .B1(n2990), .B2(n36534), .ZN(
        n9003) );
  OAI22_X1 U1744 ( .A1(n38588), .A2(n38853), .B1(n38582), .B2(n36535), .ZN(
        n9004) );
  OAI22_X1 U1745 ( .A1(n38588), .A2(n38860), .B1(n38582), .B2(n36536), .ZN(
        n9005) );
  OAI22_X1 U1746 ( .A1(n38588), .A2(n38867), .B1(n38582), .B2(n36537), .ZN(
        n9006) );
  OAI22_X1 U1747 ( .A1(n38588), .A2(n38874), .B1(n38582), .B2(n36538), .ZN(
        n9007) );
  OAI22_X1 U1748 ( .A1(n38588), .A2(n38881), .B1(n38582), .B2(n36539), .ZN(
        n9008) );
  OAI22_X1 U1749 ( .A1(n38589), .A2(n38888), .B1(n38582), .B2(n36540), .ZN(
        n9009) );
  OAI22_X1 U1750 ( .A1(n38589), .A2(n38895), .B1(n2990), .B2(n36541), .ZN(
        n9010) );
  OAI22_X1 U1751 ( .A1(n38599), .A2(n38846), .B1(n2955), .B2(n36022), .ZN(
        n9035) );
  OAI22_X1 U1752 ( .A1(n38600), .A2(n38853), .B1(n2955), .B2(n36023), .ZN(
        n9036) );
  OAI22_X1 U1753 ( .A1(n38600), .A2(n38860), .B1(n2955), .B2(n36024), .ZN(
        n9037) );
  OAI22_X1 U1754 ( .A1(n38600), .A2(n38867), .B1(n38594), .B2(n36025), .ZN(
        n9038) );
  OAI22_X1 U1755 ( .A1(n38600), .A2(n38874), .B1(n38594), .B2(n36026), .ZN(
        n9039) );
  OAI22_X1 U1756 ( .A1(n38600), .A2(n38881), .B1(n38594), .B2(n36027), .ZN(
        n9040) );
  OAI22_X1 U1757 ( .A1(n38601), .A2(n38888), .B1(n38594), .B2(n36028), .ZN(
        n9041) );
  OAI22_X1 U1758 ( .A1(n38601), .A2(n38895), .B1(n2955), .B2(n36029), .ZN(
        n9042) );
  OAI22_X1 U1759 ( .A1(n38635), .A2(n38846), .B1(n2850), .B2(n35190), .ZN(
        n9131) );
  OAI22_X1 U1760 ( .A1(n38636), .A2(n38853), .B1(n2850), .B2(n35191), .ZN(
        n9132) );
  OAI22_X1 U1761 ( .A1(n38636), .A2(n38860), .B1(n2850), .B2(n35192), .ZN(
        n9133) );
  OAI22_X1 U1762 ( .A1(n38636), .A2(n38867), .B1(n38630), .B2(n35193), .ZN(
        n9134) );
  OAI22_X1 U1763 ( .A1(n38636), .A2(n38874), .B1(n38630), .B2(n35194), .ZN(
        n9135) );
  OAI22_X1 U1764 ( .A1(n38636), .A2(n38881), .B1(n38630), .B2(n35195), .ZN(
        n9136) );
  OAI22_X1 U1765 ( .A1(n38637), .A2(n38888), .B1(n38630), .B2(n35196), .ZN(
        n9137) );
  OAI22_X1 U1766 ( .A1(n38637), .A2(n38895), .B1(n2850), .B2(n35197), .ZN(
        n9138) );
  OAI22_X1 U1767 ( .A1(n38647), .A2(n38846), .B1(n2815), .B2(n36214), .ZN(
        n9163) );
  OAI22_X1 U1768 ( .A1(n38648), .A2(n38853), .B1(n38642), .B2(n36215), .ZN(
        n9164) );
  OAI22_X1 U1769 ( .A1(n38648), .A2(n38860), .B1(n38642), .B2(n36216), .ZN(
        n9165) );
  OAI22_X1 U1770 ( .A1(n38648), .A2(n38867), .B1(n38642), .B2(n36217), .ZN(
        n9166) );
  OAI22_X1 U1771 ( .A1(n38648), .A2(n38874), .B1(n38642), .B2(n36218), .ZN(
        n9167) );
  OAI22_X1 U1772 ( .A1(n38648), .A2(n38881), .B1(n38642), .B2(n36219), .ZN(
        n9168) );
  OAI22_X1 U1773 ( .A1(n38649), .A2(n38888), .B1(n38642), .B2(n36220), .ZN(
        n9169) );
  OAI22_X1 U1774 ( .A1(n38649), .A2(n38895), .B1(n2815), .B2(n36221), .ZN(
        n9170) );
  OAI22_X1 U1775 ( .A1(n38659), .A2(n38846), .B1(n2778), .B2(n35702), .ZN(
        n9195) );
  OAI22_X1 U1776 ( .A1(n38660), .A2(n38853), .B1(n38654), .B2(n35703), .ZN(
        n9196) );
  OAI22_X1 U1777 ( .A1(n38660), .A2(n38860), .B1(n38654), .B2(n35704), .ZN(
        n9197) );
  OAI22_X1 U1778 ( .A1(n38660), .A2(n38867), .B1(n38654), .B2(n35705), .ZN(
        n9198) );
  OAI22_X1 U1779 ( .A1(n38660), .A2(n38874), .B1(n38654), .B2(n35706), .ZN(
        n9199) );
  OAI22_X1 U1780 ( .A1(n38660), .A2(n38881), .B1(n38654), .B2(n35707), .ZN(
        n9200) );
  OAI22_X1 U1781 ( .A1(n38661), .A2(n38888), .B1(n38654), .B2(n35708), .ZN(
        n9201) );
  OAI22_X1 U1782 ( .A1(n38661), .A2(n38895), .B1(n2778), .B2(n35709), .ZN(
        n9202) );
  OAI22_X1 U1783 ( .A1(n37818), .A2(n38683), .B1(n37817), .B2(n35414), .ZN(
        n6771) );
  OAI22_X1 U1784 ( .A1(n37818), .A2(n38690), .B1(n37817), .B2(n35418), .ZN(
        n6772) );
  OAI22_X1 U1785 ( .A1(n37818), .A2(n38697), .B1(n37817), .B2(n35422), .ZN(
        n6773) );
  OAI22_X1 U1786 ( .A1(n37818), .A2(n38704), .B1(n37817), .B2(n35426), .ZN(
        n6774) );
  OAI22_X1 U1787 ( .A1(n37818), .A2(n38711), .B1(n37817), .B2(n35430), .ZN(
        n6775) );
  OAI22_X1 U1788 ( .A1(n37819), .A2(n38718), .B1(n37817), .B2(n35434), .ZN(
        n6776) );
  OAI22_X1 U1789 ( .A1(n37819), .A2(n38725), .B1(n37817), .B2(n35438), .ZN(
        n6777) );
  OAI22_X1 U1790 ( .A1(n37819), .A2(n38732), .B1(n37817), .B2(n35442), .ZN(
        n6778) );
  OAI22_X1 U1791 ( .A1(n37819), .A2(n38739), .B1(n37817), .B2(n35446), .ZN(
        n6779) );
  OAI22_X1 U1792 ( .A1(n37819), .A2(n38746), .B1(n37817), .B2(n35450), .ZN(
        n6780) );
  OAI22_X1 U1793 ( .A1(n37820), .A2(n38753), .B1(n37817), .B2(n35454), .ZN(
        n6781) );
  OAI22_X1 U1794 ( .A1(n37820), .A2(n38760), .B1(n37817), .B2(n35458), .ZN(
        n6782) );
  OAI22_X1 U1795 ( .A1(n37820), .A2(n38767), .B1(n37817), .B2(n35462), .ZN(
        n6783) );
  OAI22_X1 U1796 ( .A1(n37820), .A2(n38774), .B1(n37817), .B2(n35466), .ZN(
        n6784) );
  OAI22_X1 U1797 ( .A1(n37820), .A2(n38781), .B1(n5439), .B2(n35470), .ZN(
        n6785) );
  OAI22_X1 U1798 ( .A1(n37821), .A2(n38788), .B1(n5439), .B2(n35474), .ZN(
        n6786) );
  OAI22_X1 U1799 ( .A1(n37821), .A2(n38795), .B1(n5439), .B2(n35478), .ZN(
        n6787) );
  OAI22_X1 U1800 ( .A1(n37821), .A2(n38802), .B1(n5439), .B2(n35482), .ZN(
        n6788) );
  OAI22_X1 U1801 ( .A1(n37821), .A2(n38809), .B1(n5439), .B2(n35486), .ZN(
        n6789) );
  OAI22_X1 U1802 ( .A1(n37821), .A2(n38816), .B1(n5439), .B2(n35490), .ZN(
        n6790) );
  OAI22_X1 U1803 ( .A1(n37822), .A2(n38823), .B1(n5439), .B2(n35494), .ZN(
        n6791) );
  OAI22_X1 U1804 ( .A1(n37822), .A2(n38830), .B1(n37817), .B2(n35498), .ZN(
        n6792) );
  OAI22_X1 U1805 ( .A1(n37822), .A2(n38837), .B1(n37817), .B2(n35502), .ZN(
        n6793) );
  OAI22_X1 U1806 ( .A1(n37822), .A2(n38844), .B1(n37817), .B2(n35506), .ZN(
        n6794) );
  OAI22_X1 U1807 ( .A1(n37830), .A2(n38683), .B1(n37829), .B2(n36438), .ZN(
        n6803) );
  OAI22_X1 U1808 ( .A1(n37830), .A2(n38690), .B1(n37829), .B2(n36442), .ZN(
        n6804) );
  OAI22_X1 U1809 ( .A1(n37830), .A2(n38697), .B1(n37829), .B2(n36446), .ZN(
        n6805) );
  OAI22_X1 U1810 ( .A1(n37830), .A2(n38704), .B1(n37829), .B2(n36450), .ZN(
        n6806) );
  OAI22_X1 U1811 ( .A1(n37830), .A2(n38711), .B1(n37829), .B2(n36454), .ZN(
        n6807) );
  OAI22_X1 U1812 ( .A1(n37831), .A2(n38718), .B1(n37829), .B2(n36458), .ZN(
        n6808) );
  OAI22_X1 U1813 ( .A1(n37831), .A2(n38725), .B1(n37829), .B2(n36462), .ZN(
        n6809) );
  OAI22_X1 U1814 ( .A1(n37831), .A2(n38732), .B1(n37829), .B2(n36466), .ZN(
        n6810) );
  OAI22_X1 U1815 ( .A1(n37831), .A2(n38739), .B1(n37829), .B2(n36470), .ZN(
        n6811) );
  OAI22_X1 U1816 ( .A1(n37831), .A2(n38746), .B1(n37829), .B2(n36474), .ZN(
        n6812) );
  OAI22_X1 U1817 ( .A1(n37832), .A2(n38753), .B1(n37829), .B2(n36478), .ZN(
        n6813) );
  OAI22_X1 U1818 ( .A1(n37832), .A2(n38760), .B1(n37829), .B2(n36482), .ZN(
        n6814) );
  OAI22_X1 U1819 ( .A1(n37832), .A2(n38767), .B1(n37829), .B2(n36486), .ZN(
        n6815) );
  OAI22_X1 U1820 ( .A1(n37832), .A2(n38774), .B1(n37829), .B2(n36490), .ZN(
        n6816) );
  OAI22_X1 U1821 ( .A1(n37832), .A2(n38781), .B1(n5404), .B2(n36494), .ZN(
        n6817) );
  OAI22_X1 U1822 ( .A1(n37833), .A2(n38788), .B1(n5404), .B2(n36498), .ZN(
        n6818) );
  OAI22_X1 U1823 ( .A1(n37833), .A2(n38795), .B1(n5404), .B2(n36502), .ZN(
        n6819) );
  OAI22_X1 U1824 ( .A1(n37833), .A2(n38802), .B1(n5404), .B2(n36506), .ZN(
        n6820) );
  OAI22_X1 U1825 ( .A1(n37833), .A2(n38809), .B1(n5404), .B2(n36510), .ZN(
        n6821) );
  OAI22_X1 U1826 ( .A1(n37833), .A2(n38816), .B1(n5404), .B2(n36514), .ZN(
        n6822) );
  OAI22_X1 U1827 ( .A1(n37834), .A2(n38823), .B1(n5404), .B2(n36518), .ZN(
        n6823) );
  OAI22_X1 U1828 ( .A1(n37834), .A2(n38830), .B1(n37829), .B2(n36522), .ZN(
        n6824) );
  OAI22_X1 U1829 ( .A1(n37834), .A2(n38837), .B1(n37829), .B2(n36526), .ZN(
        n6825) );
  OAI22_X1 U1830 ( .A1(n37834), .A2(n38844), .B1(n37829), .B2(n36530), .ZN(
        n6826) );
  OAI22_X1 U1831 ( .A1(n37842), .A2(n38683), .B1(n37841), .B2(n35926), .ZN(
        n6835) );
  OAI22_X1 U1832 ( .A1(n37842), .A2(n38690), .B1(n37841), .B2(n35930), .ZN(
        n6836) );
  OAI22_X1 U1833 ( .A1(n37842), .A2(n38697), .B1(n37841), .B2(n35934), .ZN(
        n6837) );
  OAI22_X1 U1834 ( .A1(n37842), .A2(n38704), .B1(n37841), .B2(n35938), .ZN(
        n6838) );
  OAI22_X1 U1835 ( .A1(n37842), .A2(n38711), .B1(n37841), .B2(n35942), .ZN(
        n6839) );
  OAI22_X1 U1836 ( .A1(n37843), .A2(n38718), .B1(n37841), .B2(n35946), .ZN(
        n6840) );
  OAI22_X1 U1837 ( .A1(n37843), .A2(n38725), .B1(n37841), .B2(n35950), .ZN(
        n6841) );
  OAI22_X1 U1838 ( .A1(n37843), .A2(n38732), .B1(n37841), .B2(n35954), .ZN(
        n6842) );
  OAI22_X1 U1839 ( .A1(n37843), .A2(n38739), .B1(n37841), .B2(n35958), .ZN(
        n6843) );
  OAI22_X1 U1840 ( .A1(n37843), .A2(n38746), .B1(n37841), .B2(n35962), .ZN(
        n6844) );
  OAI22_X1 U1841 ( .A1(n37844), .A2(n38753), .B1(n37841), .B2(n35966), .ZN(
        n6845) );
  OAI22_X1 U1842 ( .A1(n37844), .A2(n38760), .B1(n37841), .B2(n35970), .ZN(
        n6846) );
  OAI22_X1 U1843 ( .A1(n37844), .A2(n38767), .B1(n37841), .B2(n35974), .ZN(
        n6847) );
  OAI22_X1 U1844 ( .A1(n37844), .A2(n38774), .B1(n37841), .B2(n35978), .ZN(
        n6848) );
  OAI22_X1 U1845 ( .A1(n37844), .A2(n38781), .B1(n5369), .B2(n35982), .ZN(
        n6849) );
  OAI22_X1 U1846 ( .A1(n37845), .A2(n38788), .B1(n5369), .B2(n35986), .ZN(
        n6850) );
  OAI22_X1 U1847 ( .A1(n37845), .A2(n38795), .B1(n5369), .B2(n35990), .ZN(
        n6851) );
  OAI22_X1 U1848 ( .A1(n37845), .A2(n38802), .B1(n5369), .B2(n35994), .ZN(
        n6852) );
  OAI22_X1 U1849 ( .A1(n37845), .A2(n38809), .B1(n5369), .B2(n35998), .ZN(
        n6853) );
  OAI22_X1 U1850 ( .A1(n37845), .A2(n38816), .B1(n5369), .B2(n36002), .ZN(
        n6854) );
  OAI22_X1 U1851 ( .A1(n37846), .A2(n38823), .B1(n5369), .B2(n36006), .ZN(
        n6855) );
  OAI22_X1 U1852 ( .A1(n37846), .A2(n38830), .B1(n37841), .B2(n36010), .ZN(
        n6856) );
  OAI22_X1 U1853 ( .A1(n37846), .A2(n38837), .B1(n37841), .B2(n36014), .ZN(
        n6857) );
  OAI22_X1 U1854 ( .A1(n37846), .A2(n38844), .B1(n37841), .B2(n36018), .ZN(
        n6858) );
  OAI22_X1 U1855 ( .A1(n37872), .A2(n38683), .B1(n37871), .B2(n35198), .ZN(
        n6931) );
  OAI22_X1 U1856 ( .A1(n37872), .A2(n38690), .B1(n37871), .B2(n35199), .ZN(
        n6932) );
  OAI22_X1 U1857 ( .A1(n37872), .A2(n38697), .B1(n37871), .B2(n35200), .ZN(
        n6933) );
  OAI22_X1 U1858 ( .A1(n37872), .A2(n38704), .B1(n37871), .B2(n35201), .ZN(
        n6934) );
  OAI22_X1 U1859 ( .A1(n37872), .A2(n38711), .B1(n37871), .B2(n35202), .ZN(
        n6935) );
  OAI22_X1 U1860 ( .A1(n37873), .A2(n38718), .B1(n37871), .B2(n35203), .ZN(
        n6936) );
  OAI22_X1 U1861 ( .A1(n37873), .A2(n38725), .B1(n37871), .B2(n35204), .ZN(
        n6937) );
  OAI22_X1 U1862 ( .A1(n37873), .A2(n38732), .B1(n37871), .B2(n35205), .ZN(
        n6938) );
  OAI22_X1 U1863 ( .A1(n37873), .A2(n38739), .B1(n37871), .B2(n35206), .ZN(
        n6939) );
  OAI22_X1 U1864 ( .A1(n37873), .A2(n38746), .B1(n37871), .B2(n35207), .ZN(
        n6940) );
  OAI22_X1 U1865 ( .A1(n37874), .A2(n38753), .B1(n37871), .B2(n35208), .ZN(
        n6941) );
  OAI22_X1 U1866 ( .A1(n37874), .A2(n38760), .B1(n37871), .B2(n35209), .ZN(
        n6942) );
  OAI22_X1 U1867 ( .A1(n37874), .A2(n38767), .B1(n37871), .B2(n35210), .ZN(
        n6943) );
  OAI22_X1 U1868 ( .A1(n37874), .A2(n38774), .B1(n37871), .B2(n35211), .ZN(
        n6944) );
  OAI22_X1 U1869 ( .A1(n37874), .A2(n38781), .B1(n5264), .B2(n35212), .ZN(
        n6945) );
  OAI22_X1 U1870 ( .A1(n37875), .A2(n38788), .B1(n5264), .B2(n35213), .ZN(
        n6946) );
  OAI22_X1 U1871 ( .A1(n37875), .A2(n38795), .B1(n5264), .B2(n35214), .ZN(
        n6947) );
  OAI22_X1 U1872 ( .A1(n37875), .A2(n38802), .B1(n5264), .B2(n35215), .ZN(
        n6948) );
  OAI22_X1 U1873 ( .A1(n37875), .A2(n38809), .B1(n5264), .B2(n35216), .ZN(
        n6949) );
  OAI22_X1 U1874 ( .A1(n37875), .A2(n38816), .B1(n5264), .B2(n35217), .ZN(
        n6950) );
  OAI22_X1 U1875 ( .A1(n37876), .A2(n38823), .B1(n5264), .B2(n35218), .ZN(
        n6951) );
  OAI22_X1 U1876 ( .A1(n37876), .A2(n38830), .B1(n37871), .B2(n35219), .ZN(
        n6952) );
  OAI22_X1 U1877 ( .A1(n37876), .A2(n38837), .B1(n37871), .B2(n35220), .ZN(
        n6953) );
  OAI22_X1 U1878 ( .A1(n37876), .A2(n38844), .B1(n37871), .B2(n35221), .ZN(
        n6954) );
  OAI22_X1 U1879 ( .A1(n37884), .A2(n38683), .B1(n37883), .B2(n36222), .ZN(
        n6963) );
  OAI22_X1 U1880 ( .A1(n37884), .A2(n38690), .B1(n37883), .B2(n36223), .ZN(
        n6964) );
  OAI22_X1 U1881 ( .A1(n37884), .A2(n38697), .B1(n37883), .B2(n36224), .ZN(
        n6965) );
  OAI22_X1 U1882 ( .A1(n37884), .A2(n38704), .B1(n37883), .B2(n36225), .ZN(
        n6966) );
  OAI22_X1 U1883 ( .A1(n37884), .A2(n38711), .B1(n37883), .B2(n36226), .ZN(
        n6967) );
  OAI22_X1 U1884 ( .A1(n37885), .A2(n38718), .B1(n37883), .B2(n36227), .ZN(
        n6968) );
  OAI22_X1 U1885 ( .A1(n37885), .A2(n38725), .B1(n37883), .B2(n36228), .ZN(
        n6969) );
  OAI22_X1 U1886 ( .A1(n37885), .A2(n38732), .B1(n37883), .B2(n36229), .ZN(
        n6970) );
  OAI22_X1 U1887 ( .A1(n37885), .A2(n38739), .B1(n37883), .B2(n36230), .ZN(
        n6971) );
  OAI22_X1 U1888 ( .A1(n37885), .A2(n38746), .B1(n37883), .B2(n36231), .ZN(
        n6972) );
  OAI22_X1 U1889 ( .A1(n37886), .A2(n38753), .B1(n37883), .B2(n36232), .ZN(
        n6973) );
  OAI22_X1 U1890 ( .A1(n37886), .A2(n38760), .B1(n37883), .B2(n36233), .ZN(
        n6974) );
  OAI22_X1 U1891 ( .A1(n37886), .A2(n38767), .B1(n37883), .B2(n36234), .ZN(
        n6975) );
  OAI22_X1 U1892 ( .A1(n37886), .A2(n38774), .B1(n37883), .B2(n36235), .ZN(
        n6976) );
  OAI22_X1 U1893 ( .A1(n37886), .A2(n38781), .B1(n5229), .B2(n36236), .ZN(
        n6977) );
  OAI22_X1 U1894 ( .A1(n37887), .A2(n38788), .B1(n5229), .B2(n36237), .ZN(
        n6978) );
  OAI22_X1 U1895 ( .A1(n37887), .A2(n38795), .B1(n5229), .B2(n36238), .ZN(
        n6979) );
  OAI22_X1 U1896 ( .A1(n37887), .A2(n38802), .B1(n5229), .B2(n36239), .ZN(
        n6980) );
  OAI22_X1 U1897 ( .A1(n37887), .A2(n38809), .B1(n5229), .B2(n36240), .ZN(
        n6981) );
  OAI22_X1 U1898 ( .A1(n37887), .A2(n38816), .B1(n5229), .B2(n36241), .ZN(
        n6982) );
  OAI22_X1 U1899 ( .A1(n37888), .A2(n38823), .B1(n5229), .B2(n36242), .ZN(
        n6983) );
  OAI22_X1 U1900 ( .A1(n37888), .A2(n38830), .B1(n37883), .B2(n36243), .ZN(
        n6984) );
  OAI22_X1 U1901 ( .A1(n37888), .A2(n38837), .B1(n37883), .B2(n36244), .ZN(
        n6985) );
  OAI22_X1 U1902 ( .A1(n37888), .A2(n38844), .B1(n37883), .B2(n36245), .ZN(
        n6986) );
  OAI22_X1 U1903 ( .A1(n37896), .A2(n38683), .B1(n37895), .B2(n35710), .ZN(
        n6995) );
  OAI22_X1 U1904 ( .A1(n37896), .A2(n38690), .B1(n37895), .B2(n35711), .ZN(
        n6996) );
  OAI22_X1 U1905 ( .A1(n37896), .A2(n38697), .B1(n37895), .B2(n35712), .ZN(
        n6997) );
  OAI22_X1 U1906 ( .A1(n37896), .A2(n38704), .B1(n37895), .B2(n35713), .ZN(
        n6998) );
  OAI22_X1 U1907 ( .A1(n37896), .A2(n38711), .B1(n37895), .B2(n35714), .ZN(
        n6999) );
  OAI22_X1 U1908 ( .A1(n37897), .A2(n38718), .B1(n37895), .B2(n35715), .ZN(
        n7000) );
  OAI22_X1 U1909 ( .A1(n37897), .A2(n38725), .B1(n37895), .B2(n35716), .ZN(
        n7001) );
  OAI22_X1 U1910 ( .A1(n37897), .A2(n38732), .B1(n37895), .B2(n35717), .ZN(
        n7002) );
  OAI22_X1 U1911 ( .A1(n37897), .A2(n38739), .B1(n37895), .B2(n35718), .ZN(
        n7003) );
  OAI22_X1 U1912 ( .A1(n37897), .A2(n38746), .B1(n37895), .B2(n35719), .ZN(
        n7004) );
  OAI22_X1 U1913 ( .A1(n37898), .A2(n38753), .B1(n37895), .B2(n35720), .ZN(
        n7005) );
  OAI22_X1 U1914 ( .A1(n37898), .A2(n38760), .B1(n37895), .B2(n35721), .ZN(
        n7006) );
  OAI22_X1 U1915 ( .A1(n37898), .A2(n38767), .B1(n37895), .B2(n35722), .ZN(
        n7007) );
  OAI22_X1 U1916 ( .A1(n37898), .A2(n38774), .B1(n37895), .B2(n35723), .ZN(
        n7008) );
  OAI22_X1 U1917 ( .A1(n37898), .A2(n38781), .B1(n5194), .B2(n35724), .ZN(
        n7009) );
  OAI22_X1 U1918 ( .A1(n37899), .A2(n38788), .B1(n5194), .B2(n35725), .ZN(
        n7010) );
  OAI22_X1 U1919 ( .A1(n37899), .A2(n38795), .B1(n5194), .B2(n35726), .ZN(
        n7011) );
  OAI22_X1 U1920 ( .A1(n37899), .A2(n38802), .B1(n5194), .B2(n35727), .ZN(
        n7012) );
  OAI22_X1 U1921 ( .A1(n37899), .A2(n38809), .B1(n5194), .B2(n35728), .ZN(
        n7013) );
  OAI22_X1 U1922 ( .A1(n37899), .A2(n38816), .B1(n5194), .B2(n35729), .ZN(
        n7014) );
  OAI22_X1 U1923 ( .A1(n37900), .A2(n38823), .B1(n5194), .B2(n35730), .ZN(
        n7015) );
  OAI22_X1 U1924 ( .A1(n37900), .A2(n38830), .B1(n37895), .B2(n35731), .ZN(
        n7016) );
  OAI22_X1 U1925 ( .A1(n37900), .A2(n38837), .B1(n37895), .B2(n35732), .ZN(
        n7017) );
  OAI22_X1 U1926 ( .A1(n37900), .A2(n38844), .B1(n37895), .B2(n35733), .ZN(
        n7018) );
  OAI22_X1 U1927 ( .A1(n37926), .A2(n38683), .B1(n37925), .B2(n35222), .ZN(
        n7091) );
  OAI22_X1 U1928 ( .A1(n37926), .A2(n38690), .B1(n37925), .B2(n35223), .ZN(
        n7092) );
  OAI22_X1 U1929 ( .A1(n37926), .A2(n38697), .B1(n37925), .B2(n35224), .ZN(
        n7093) );
  OAI22_X1 U1930 ( .A1(n37926), .A2(n38704), .B1(n37925), .B2(n35225), .ZN(
        n7094) );
  OAI22_X1 U1931 ( .A1(n37926), .A2(n38711), .B1(n37925), .B2(n35226), .ZN(
        n7095) );
  OAI22_X1 U1932 ( .A1(n37927), .A2(n38718), .B1(n37925), .B2(n35227), .ZN(
        n7096) );
  OAI22_X1 U1933 ( .A1(n37927), .A2(n38725), .B1(n37925), .B2(n35228), .ZN(
        n7097) );
  OAI22_X1 U1934 ( .A1(n37927), .A2(n38732), .B1(n37925), .B2(n35229), .ZN(
        n7098) );
  OAI22_X1 U1935 ( .A1(n37927), .A2(n38739), .B1(n37925), .B2(n35230), .ZN(
        n7099) );
  OAI22_X1 U1936 ( .A1(n37927), .A2(n38746), .B1(n37925), .B2(n35231), .ZN(
        n7100) );
  OAI22_X1 U1937 ( .A1(n37928), .A2(n38753), .B1(n37925), .B2(n35232), .ZN(
        n7101) );
  OAI22_X1 U1938 ( .A1(n37928), .A2(n38760), .B1(n37925), .B2(n35233), .ZN(
        n7102) );
  OAI22_X1 U1939 ( .A1(n37928), .A2(n38767), .B1(n37925), .B2(n35234), .ZN(
        n7103) );
  OAI22_X1 U1940 ( .A1(n37928), .A2(n38774), .B1(n37925), .B2(n35235), .ZN(
        n7104) );
  OAI22_X1 U1941 ( .A1(n37928), .A2(n38781), .B1(n5089), .B2(n35236), .ZN(
        n7105) );
  OAI22_X1 U1942 ( .A1(n37929), .A2(n38788), .B1(n5089), .B2(n35237), .ZN(
        n7106) );
  OAI22_X1 U1943 ( .A1(n37929), .A2(n38795), .B1(n5089), .B2(n35238), .ZN(
        n7107) );
  OAI22_X1 U1944 ( .A1(n37929), .A2(n38802), .B1(n5089), .B2(n35239), .ZN(
        n7108) );
  OAI22_X1 U1945 ( .A1(n37929), .A2(n38809), .B1(n5089), .B2(n35240), .ZN(
        n7109) );
  OAI22_X1 U1946 ( .A1(n37929), .A2(n38816), .B1(n5089), .B2(n35241), .ZN(
        n7110) );
  OAI22_X1 U1947 ( .A1(n37930), .A2(n38823), .B1(n5089), .B2(n35242), .ZN(
        n7111) );
  OAI22_X1 U1948 ( .A1(n37930), .A2(n38830), .B1(n37925), .B2(n35243), .ZN(
        n7112) );
  OAI22_X1 U1949 ( .A1(n37930), .A2(n38837), .B1(n37925), .B2(n35244), .ZN(
        n7113) );
  OAI22_X1 U1950 ( .A1(n37930), .A2(n38844), .B1(n37925), .B2(n35245), .ZN(
        n7114) );
  OAI22_X1 U1951 ( .A1(n37938), .A2(n38682), .B1(n37937), .B2(n36246), .ZN(
        n7123) );
  OAI22_X1 U1952 ( .A1(n37938), .A2(n38689), .B1(n37937), .B2(n36247), .ZN(
        n7124) );
  OAI22_X1 U1953 ( .A1(n37938), .A2(n38696), .B1(n37937), .B2(n36248), .ZN(
        n7125) );
  OAI22_X1 U1954 ( .A1(n37938), .A2(n38703), .B1(n37937), .B2(n36249), .ZN(
        n7126) );
  OAI22_X1 U1955 ( .A1(n37938), .A2(n38710), .B1(n37937), .B2(n36250), .ZN(
        n7127) );
  OAI22_X1 U1956 ( .A1(n37939), .A2(n38717), .B1(n37937), .B2(n36251), .ZN(
        n7128) );
  OAI22_X1 U1957 ( .A1(n37939), .A2(n38724), .B1(n37937), .B2(n36252), .ZN(
        n7129) );
  OAI22_X1 U1958 ( .A1(n37939), .A2(n38731), .B1(n37937), .B2(n36253), .ZN(
        n7130) );
  OAI22_X1 U1959 ( .A1(n37939), .A2(n38738), .B1(n37937), .B2(n36254), .ZN(
        n7131) );
  OAI22_X1 U1960 ( .A1(n37939), .A2(n38745), .B1(n37937), .B2(n36255), .ZN(
        n7132) );
  OAI22_X1 U1961 ( .A1(n37940), .A2(n38752), .B1(n37937), .B2(n36256), .ZN(
        n7133) );
  OAI22_X1 U1962 ( .A1(n37940), .A2(n38759), .B1(n37937), .B2(n36257), .ZN(
        n7134) );
  OAI22_X1 U1963 ( .A1(n37940), .A2(n38766), .B1(n37937), .B2(n36258), .ZN(
        n7135) );
  OAI22_X1 U1964 ( .A1(n37940), .A2(n38773), .B1(n37937), .B2(n36259), .ZN(
        n7136) );
  OAI22_X1 U1965 ( .A1(n37940), .A2(n38780), .B1(n5054), .B2(n36260), .ZN(
        n7137) );
  OAI22_X1 U1966 ( .A1(n37941), .A2(n38787), .B1(n5054), .B2(n36261), .ZN(
        n7138) );
  OAI22_X1 U1967 ( .A1(n37941), .A2(n38794), .B1(n5054), .B2(n36262), .ZN(
        n7139) );
  OAI22_X1 U1968 ( .A1(n37941), .A2(n38801), .B1(n5054), .B2(n36263), .ZN(
        n7140) );
  OAI22_X1 U1969 ( .A1(n37941), .A2(n38808), .B1(n5054), .B2(n36264), .ZN(
        n7141) );
  OAI22_X1 U1970 ( .A1(n37941), .A2(n38815), .B1(n5054), .B2(n36265), .ZN(
        n7142) );
  OAI22_X1 U1971 ( .A1(n37942), .A2(n38822), .B1(n5054), .B2(n36266), .ZN(
        n7143) );
  OAI22_X1 U1972 ( .A1(n37942), .A2(n38829), .B1(n37937), .B2(n36267), .ZN(
        n7144) );
  OAI22_X1 U1973 ( .A1(n37942), .A2(n38836), .B1(n37937), .B2(n36268), .ZN(
        n7145) );
  OAI22_X1 U1974 ( .A1(n37942), .A2(n38843), .B1(n37937), .B2(n36269), .ZN(
        n7146) );
  OAI22_X1 U1975 ( .A1(n37950), .A2(n38682), .B1(n37949), .B2(n35734), .ZN(
        n7155) );
  OAI22_X1 U1976 ( .A1(n37950), .A2(n38689), .B1(n37949), .B2(n35735), .ZN(
        n7156) );
  OAI22_X1 U1977 ( .A1(n37950), .A2(n38696), .B1(n37949), .B2(n35736), .ZN(
        n7157) );
  OAI22_X1 U1978 ( .A1(n37950), .A2(n38703), .B1(n37949), .B2(n35737), .ZN(
        n7158) );
  OAI22_X1 U1979 ( .A1(n37950), .A2(n38710), .B1(n37949), .B2(n35738), .ZN(
        n7159) );
  OAI22_X1 U1980 ( .A1(n37951), .A2(n38717), .B1(n37949), .B2(n35739), .ZN(
        n7160) );
  OAI22_X1 U1981 ( .A1(n37951), .A2(n38724), .B1(n37949), .B2(n35740), .ZN(
        n7161) );
  OAI22_X1 U1982 ( .A1(n37951), .A2(n38731), .B1(n37949), .B2(n35741), .ZN(
        n7162) );
  OAI22_X1 U1983 ( .A1(n37951), .A2(n38738), .B1(n37949), .B2(n35742), .ZN(
        n7163) );
  OAI22_X1 U1984 ( .A1(n37951), .A2(n38745), .B1(n37949), .B2(n35743), .ZN(
        n7164) );
  OAI22_X1 U1985 ( .A1(n37952), .A2(n38752), .B1(n37949), .B2(n35744), .ZN(
        n7165) );
  OAI22_X1 U1986 ( .A1(n37952), .A2(n38759), .B1(n37949), .B2(n35745), .ZN(
        n7166) );
  OAI22_X1 U1987 ( .A1(n37952), .A2(n38766), .B1(n37949), .B2(n35746), .ZN(
        n7167) );
  OAI22_X1 U1988 ( .A1(n37952), .A2(n38773), .B1(n37949), .B2(n35747), .ZN(
        n7168) );
  OAI22_X1 U1989 ( .A1(n37952), .A2(n38780), .B1(n5019), .B2(n35748), .ZN(
        n7169) );
  OAI22_X1 U1990 ( .A1(n37953), .A2(n38787), .B1(n5019), .B2(n35749), .ZN(
        n7170) );
  OAI22_X1 U1991 ( .A1(n37953), .A2(n38794), .B1(n5019), .B2(n35750), .ZN(
        n7171) );
  OAI22_X1 U1992 ( .A1(n37953), .A2(n38801), .B1(n5019), .B2(n35751), .ZN(
        n7172) );
  OAI22_X1 U1993 ( .A1(n37953), .A2(n38808), .B1(n5019), .B2(n35752), .ZN(
        n7173) );
  OAI22_X1 U1994 ( .A1(n37953), .A2(n38815), .B1(n5019), .B2(n35753), .ZN(
        n7174) );
  OAI22_X1 U1995 ( .A1(n37954), .A2(n38822), .B1(n5019), .B2(n35754), .ZN(
        n7175) );
  OAI22_X1 U1996 ( .A1(n37954), .A2(n38829), .B1(n37949), .B2(n35755), .ZN(
        n7176) );
  OAI22_X1 U1997 ( .A1(n37954), .A2(n38836), .B1(n37949), .B2(n35756), .ZN(
        n7177) );
  OAI22_X1 U1998 ( .A1(n37954), .A2(n38843), .B1(n37949), .B2(n35757), .ZN(
        n7178) );
  OAI22_X1 U1999 ( .A1(n37971), .A2(n38682), .B1(n37970), .B2(n36078), .ZN(
        n7219) );
  OAI22_X1 U2000 ( .A1(n37971), .A2(n38689), .B1(n37970), .B2(n36080), .ZN(
        n7220) );
  OAI22_X1 U2001 ( .A1(n37971), .A2(n38696), .B1(n37970), .B2(n36082), .ZN(
        n7221) );
  OAI22_X1 U2002 ( .A1(n37971), .A2(n38703), .B1(n37970), .B2(n36084), .ZN(
        n7222) );
  OAI22_X1 U2003 ( .A1(n37971), .A2(n38710), .B1(n37970), .B2(n36086), .ZN(
        n7223) );
  OAI22_X1 U2004 ( .A1(n37972), .A2(n38717), .B1(n37970), .B2(n36088), .ZN(
        n7224) );
  OAI22_X1 U2005 ( .A1(n37972), .A2(n38724), .B1(n37970), .B2(n36090), .ZN(
        n7225) );
  OAI22_X1 U2006 ( .A1(n37972), .A2(n38731), .B1(n37970), .B2(n36092), .ZN(
        n7226) );
  OAI22_X1 U2007 ( .A1(n37972), .A2(n38738), .B1(n37970), .B2(n36094), .ZN(
        n7227) );
  OAI22_X1 U2008 ( .A1(n37972), .A2(n38745), .B1(n37970), .B2(n36096), .ZN(
        n7228) );
  OAI22_X1 U2009 ( .A1(n37973), .A2(n38752), .B1(n37970), .B2(n36098), .ZN(
        n7229) );
  OAI22_X1 U2010 ( .A1(n37973), .A2(n38759), .B1(n37970), .B2(n36100), .ZN(
        n7230) );
  OAI22_X1 U2011 ( .A1(n37973), .A2(n38766), .B1(n37970), .B2(n36102), .ZN(
        n7231) );
  OAI22_X1 U2012 ( .A1(n37973), .A2(n38773), .B1(n37970), .B2(n36104), .ZN(
        n7232) );
  OAI22_X1 U2013 ( .A1(n37973), .A2(n38780), .B1(n4948), .B2(n36106), .ZN(
        n7233) );
  OAI22_X1 U2014 ( .A1(n37974), .A2(n38787), .B1(n4948), .B2(n36108), .ZN(
        n7234) );
  OAI22_X1 U2015 ( .A1(n37974), .A2(n38794), .B1(n4948), .B2(n36110), .ZN(
        n7235) );
  OAI22_X1 U2016 ( .A1(n37974), .A2(n38801), .B1(n4948), .B2(n36112), .ZN(
        n7236) );
  OAI22_X1 U2017 ( .A1(n37974), .A2(n38808), .B1(n4948), .B2(n36114), .ZN(
        n7237) );
  OAI22_X1 U2018 ( .A1(n37974), .A2(n38815), .B1(n4948), .B2(n36116), .ZN(
        n7238) );
  OAI22_X1 U2019 ( .A1(n37975), .A2(n38822), .B1(n4948), .B2(n36118), .ZN(
        n7239) );
  OAI22_X1 U2020 ( .A1(n37975), .A2(n38829), .B1(n37970), .B2(n36120), .ZN(
        n7240) );
  OAI22_X1 U2021 ( .A1(n37975), .A2(n38836), .B1(n37970), .B2(n36122), .ZN(
        n7241) );
  OAI22_X1 U2022 ( .A1(n37975), .A2(n38843), .B1(n37970), .B2(n36124), .ZN(
        n7242) );
  OAI22_X1 U2023 ( .A1(n37983), .A2(n38682), .B1(n37982), .B2(n35614), .ZN(
        n7251) );
  OAI22_X1 U2024 ( .A1(n37983), .A2(n38689), .B1(n37982), .B2(n35616), .ZN(
        n7252) );
  OAI22_X1 U2025 ( .A1(n37983), .A2(n38696), .B1(n37982), .B2(n35618), .ZN(
        n7253) );
  OAI22_X1 U2026 ( .A1(n37983), .A2(n38703), .B1(n37982), .B2(n35620), .ZN(
        n7254) );
  OAI22_X1 U2027 ( .A1(n37983), .A2(n38710), .B1(n37982), .B2(n35622), .ZN(
        n7255) );
  OAI22_X1 U2028 ( .A1(n37984), .A2(n38717), .B1(n37982), .B2(n35624), .ZN(
        n7256) );
  OAI22_X1 U2029 ( .A1(n37984), .A2(n38724), .B1(n37982), .B2(n35626), .ZN(
        n7257) );
  OAI22_X1 U2030 ( .A1(n37984), .A2(n38731), .B1(n37982), .B2(n35628), .ZN(
        n7258) );
  OAI22_X1 U2031 ( .A1(n37984), .A2(n38738), .B1(n37982), .B2(n35630), .ZN(
        n7259) );
  OAI22_X1 U2032 ( .A1(n37984), .A2(n38745), .B1(n37982), .B2(n35632), .ZN(
        n7260) );
  OAI22_X1 U2033 ( .A1(n37985), .A2(n38752), .B1(n37982), .B2(n35634), .ZN(
        n7261) );
  OAI22_X1 U2034 ( .A1(n37985), .A2(n38759), .B1(n37982), .B2(n35636), .ZN(
        n7262) );
  OAI22_X1 U2035 ( .A1(n37985), .A2(n38766), .B1(n37982), .B2(n35638), .ZN(
        n7263) );
  OAI22_X1 U2036 ( .A1(n37985), .A2(n38773), .B1(n37982), .B2(n35640), .ZN(
        n7264) );
  OAI22_X1 U2037 ( .A1(n37985), .A2(n38780), .B1(n4913), .B2(n35642), .ZN(
        n7265) );
  OAI22_X1 U2038 ( .A1(n37986), .A2(n38787), .B1(n4913), .B2(n35644), .ZN(
        n7266) );
  OAI22_X1 U2039 ( .A1(n37986), .A2(n38794), .B1(n4913), .B2(n35646), .ZN(
        n7267) );
  OAI22_X1 U2040 ( .A1(n37986), .A2(n38801), .B1(n4913), .B2(n35648), .ZN(
        n7268) );
  OAI22_X1 U2041 ( .A1(n37986), .A2(n38808), .B1(n4913), .B2(n35650), .ZN(
        n7269) );
  OAI22_X1 U2042 ( .A1(n37986), .A2(n38815), .B1(n4913), .B2(n35652), .ZN(
        n7270) );
  OAI22_X1 U2043 ( .A1(n37987), .A2(n38822), .B1(n4913), .B2(n35654), .ZN(
        n7271) );
  OAI22_X1 U2044 ( .A1(n37987), .A2(n38829), .B1(n37982), .B2(n35656), .ZN(
        n7272) );
  OAI22_X1 U2045 ( .A1(n37987), .A2(n38836), .B1(n37982), .B2(n35658), .ZN(
        n7273) );
  OAI22_X1 U2046 ( .A1(n37987), .A2(n38843), .B1(n37982), .B2(n35660), .ZN(
        n7274) );
  OAI22_X1 U2047 ( .A1(n38004), .A2(n38682), .B1(n38003), .B2(n36440), .ZN(
        n7315) );
  OAI22_X1 U2048 ( .A1(n38004), .A2(n38689), .B1(n38003), .B2(n36444), .ZN(
        n7316) );
  OAI22_X1 U2049 ( .A1(n38004), .A2(n38696), .B1(n38003), .B2(n36448), .ZN(
        n7317) );
  OAI22_X1 U2050 ( .A1(n38004), .A2(n38703), .B1(n38003), .B2(n36452), .ZN(
        n7318) );
  OAI22_X1 U2051 ( .A1(n38004), .A2(n38710), .B1(n38003), .B2(n36456), .ZN(
        n7319) );
  OAI22_X1 U2052 ( .A1(n38005), .A2(n38717), .B1(n38003), .B2(n36460), .ZN(
        n7320) );
  OAI22_X1 U2053 ( .A1(n38005), .A2(n38724), .B1(n38003), .B2(n36464), .ZN(
        n7321) );
  OAI22_X1 U2054 ( .A1(n38005), .A2(n38731), .B1(n38003), .B2(n36468), .ZN(
        n7322) );
  OAI22_X1 U2055 ( .A1(n38005), .A2(n38738), .B1(n38003), .B2(n36472), .ZN(
        n7323) );
  OAI22_X1 U2056 ( .A1(n38005), .A2(n38745), .B1(n38003), .B2(n36476), .ZN(
        n7324) );
  OAI22_X1 U2057 ( .A1(n38006), .A2(n38752), .B1(n38003), .B2(n36480), .ZN(
        n7325) );
  OAI22_X1 U2058 ( .A1(n38006), .A2(n38759), .B1(n38003), .B2(n36484), .ZN(
        n7326) );
  OAI22_X1 U2059 ( .A1(n38006), .A2(n38766), .B1(n38003), .B2(n36488), .ZN(
        n7327) );
  OAI22_X1 U2060 ( .A1(n38006), .A2(n38773), .B1(n38003), .B2(n36492), .ZN(
        n7328) );
  OAI22_X1 U2061 ( .A1(n38006), .A2(n38780), .B1(n4843), .B2(n36496), .ZN(
        n7329) );
  OAI22_X1 U2062 ( .A1(n38007), .A2(n38787), .B1(n4843), .B2(n36500), .ZN(
        n7330) );
  OAI22_X1 U2063 ( .A1(n38007), .A2(n38794), .B1(n4843), .B2(n36504), .ZN(
        n7331) );
  OAI22_X1 U2064 ( .A1(n38007), .A2(n38801), .B1(n4843), .B2(n36508), .ZN(
        n7332) );
  OAI22_X1 U2065 ( .A1(n38007), .A2(n38808), .B1(n4843), .B2(n36512), .ZN(
        n7333) );
  OAI22_X1 U2066 ( .A1(n38007), .A2(n38815), .B1(n4843), .B2(n36516), .ZN(
        n7334) );
  OAI22_X1 U2067 ( .A1(n38008), .A2(n38822), .B1(n4843), .B2(n36520), .ZN(
        n7335) );
  OAI22_X1 U2068 ( .A1(n38008), .A2(n38829), .B1(n38003), .B2(n36524), .ZN(
        n7336) );
  OAI22_X1 U2069 ( .A1(n38008), .A2(n38836), .B1(n38003), .B2(n36528), .ZN(
        n7337) );
  OAI22_X1 U2070 ( .A1(n38008), .A2(n38843), .B1(n38003), .B2(n36532), .ZN(
        n7338) );
  OAI22_X1 U2071 ( .A1(n38025), .A2(n38682), .B1(n38024), .B2(n36030), .ZN(
        n7379) );
  OAI22_X1 U2072 ( .A1(n38025), .A2(n38689), .B1(n38024), .B2(n36032), .ZN(
        n7380) );
  OAI22_X1 U2073 ( .A1(n38025), .A2(n38696), .B1(n38024), .B2(n36034), .ZN(
        n7381) );
  OAI22_X1 U2074 ( .A1(n38025), .A2(n38703), .B1(n38024), .B2(n36036), .ZN(
        n7382) );
  OAI22_X1 U2075 ( .A1(n38025), .A2(n38710), .B1(n38024), .B2(n36038), .ZN(
        n7383) );
  OAI22_X1 U2076 ( .A1(n38026), .A2(n38717), .B1(n38024), .B2(n36040), .ZN(
        n7384) );
  OAI22_X1 U2077 ( .A1(n38026), .A2(n38724), .B1(n38024), .B2(n36042), .ZN(
        n7385) );
  OAI22_X1 U2078 ( .A1(n38026), .A2(n38731), .B1(n38024), .B2(n36044), .ZN(
        n7386) );
  OAI22_X1 U2079 ( .A1(n38026), .A2(n38738), .B1(n38024), .B2(n36046), .ZN(
        n7387) );
  OAI22_X1 U2080 ( .A1(n38026), .A2(n38745), .B1(n38024), .B2(n36048), .ZN(
        n7388) );
  OAI22_X1 U2081 ( .A1(n38027), .A2(n38752), .B1(n38024), .B2(n36050), .ZN(
        n7389) );
  OAI22_X1 U2082 ( .A1(n38027), .A2(n38759), .B1(n38024), .B2(n36052), .ZN(
        n7390) );
  OAI22_X1 U2083 ( .A1(n38027), .A2(n38766), .B1(n38024), .B2(n36054), .ZN(
        n7391) );
  OAI22_X1 U2084 ( .A1(n38027), .A2(n38773), .B1(n38024), .B2(n36056), .ZN(
        n7392) );
  OAI22_X1 U2085 ( .A1(n38027), .A2(n38780), .B1(n4773), .B2(n36058), .ZN(
        n7393) );
  OAI22_X1 U2086 ( .A1(n38028), .A2(n38787), .B1(n4773), .B2(n36060), .ZN(
        n7394) );
  OAI22_X1 U2087 ( .A1(n38028), .A2(n38794), .B1(n4773), .B2(n36062), .ZN(
        n7395) );
  OAI22_X1 U2088 ( .A1(n38028), .A2(n38801), .B1(n4773), .B2(n36064), .ZN(
        n7396) );
  OAI22_X1 U2089 ( .A1(n38028), .A2(n38808), .B1(n4773), .B2(n36066), .ZN(
        n7397) );
  OAI22_X1 U2090 ( .A1(n38028), .A2(n38815), .B1(n4773), .B2(n36068), .ZN(
        n7398) );
  OAI22_X1 U2091 ( .A1(n38029), .A2(n38822), .B1(n4773), .B2(n36070), .ZN(
        n7399) );
  OAI22_X1 U2092 ( .A1(n38029), .A2(n38829), .B1(n38024), .B2(n36072), .ZN(
        n7400) );
  OAI22_X1 U2093 ( .A1(n38029), .A2(n38836), .B1(n38024), .B2(n36074), .ZN(
        n7401) );
  OAI22_X1 U2094 ( .A1(n38029), .A2(n38843), .B1(n38024), .B2(n36076), .ZN(
        n7402) );
  OAI22_X1 U2095 ( .A1(n38037), .A2(n38682), .B1(n38036), .B2(n35567), .ZN(
        n7411) );
  OAI22_X1 U2096 ( .A1(n38037), .A2(n38689), .B1(n38036), .B2(n35569), .ZN(
        n7412) );
  OAI22_X1 U2097 ( .A1(n38037), .A2(n38696), .B1(n38036), .B2(n35571), .ZN(
        n7413) );
  OAI22_X1 U2098 ( .A1(n38037), .A2(n38703), .B1(n38036), .B2(n35573), .ZN(
        n7414) );
  OAI22_X1 U2099 ( .A1(n38037), .A2(n38710), .B1(n38036), .B2(n35575), .ZN(
        n7415) );
  OAI22_X1 U2100 ( .A1(n38038), .A2(n38717), .B1(n38036), .B2(n35577), .ZN(
        n7416) );
  OAI22_X1 U2101 ( .A1(n38038), .A2(n38724), .B1(n38036), .B2(n35579), .ZN(
        n7417) );
  OAI22_X1 U2102 ( .A1(n38038), .A2(n38731), .B1(n38036), .B2(n35581), .ZN(
        n7418) );
  OAI22_X1 U2103 ( .A1(n38038), .A2(n38738), .B1(n38036), .B2(n35583), .ZN(
        n7419) );
  OAI22_X1 U2104 ( .A1(n38038), .A2(n38745), .B1(n38036), .B2(n35585), .ZN(
        n7420) );
  OAI22_X1 U2105 ( .A1(n38039), .A2(n38752), .B1(n38036), .B2(n35587), .ZN(
        n7421) );
  OAI22_X1 U2106 ( .A1(n38039), .A2(n38759), .B1(n38036), .B2(n35589), .ZN(
        n7422) );
  OAI22_X1 U2107 ( .A1(n38039), .A2(n38766), .B1(n38036), .B2(n35591), .ZN(
        n7423) );
  OAI22_X1 U2108 ( .A1(n38039), .A2(n38773), .B1(n38036), .B2(n35593), .ZN(
        n7424) );
  OAI22_X1 U2109 ( .A1(n38039), .A2(n38780), .B1(n4738), .B2(n35595), .ZN(
        n7425) );
  OAI22_X1 U2110 ( .A1(n38040), .A2(n38787), .B1(n4738), .B2(n35597), .ZN(
        n7426) );
  OAI22_X1 U2111 ( .A1(n38040), .A2(n38794), .B1(n4738), .B2(n35599), .ZN(
        n7427) );
  OAI22_X1 U2112 ( .A1(n38040), .A2(n38801), .B1(n4738), .B2(n35601), .ZN(
        n7428) );
  OAI22_X1 U2113 ( .A1(n38040), .A2(n38808), .B1(n4738), .B2(n35603), .ZN(
        n7429) );
  OAI22_X1 U2114 ( .A1(n38040), .A2(n38815), .B1(n4738), .B2(n35605), .ZN(
        n7430) );
  OAI22_X1 U2115 ( .A1(n38041), .A2(n38822), .B1(n4738), .B2(n35607), .ZN(
        n7431) );
  OAI22_X1 U2116 ( .A1(n38041), .A2(n38829), .B1(n38036), .B2(n35609), .ZN(
        n7432) );
  OAI22_X1 U2117 ( .A1(n38041), .A2(n38836), .B1(n38036), .B2(n35611), .ZN(
        n7433) );
  OAI22_X1 U2118 ( .A1(n38041), .A2(n38843), .B1(n38036), .B2(n35613), .ZN(
        n7434) );
  OAI22_X1 U2119 ( .A1(n38058), .A2(n38682), .B1(n38057), .B2(n36639), .ZN(
        n7475) );
  OAI22_X1 U2120 ( .A1(n38058), .A2(n38689), .B1(n38057), .B2(n36641), .ZN(
        n7476) );
  OAI22_X1 U2121 ( .A1(n38058), .A2(n38696), .B1(n38057), .B2(n36643), .ZN(
        n7477) );
  OAI22_X1 U2122 ( .A1(n38058), .A2(n38703), .B1(n38057), .B2(n36645), .ZN(
        n7478) );
  OAI22_X1 U2123 ( .A1(n38058), .A2(n38710), .B1(n38057), .B2(n36647), .ZN(
        n7479) );
  OAI22_X1 U2124 ( .A1(n38059), .A2(n38717), .B1(n38057), .B2(n36649), .ZN(
        n7480) );
  OAI22_X1 U2125 ( .A1(n38059), .A2(n38724), .B1(n38057), .B2(n36651), .ZN(
        n7481) );
  OAI22_X1 U2126 ( .A1(n38059), .A2(n38731), .B1(n38057), .B2(n36653), .ZN(
        n7482) );
  OAI22_X1 U2127 ( .A1(n38059), .A2(n38738), .B1(n38057), .B2(n36655), .ZN(
        n7483) );
  OAI22_X1 U2128 ( .A1(n38059), .A2(n38745), .B1(n38057), .B2(n36657), .ZN(
        n7484) );
  OAI22_X1 U2129 ( .A1(n38060), .A2(n38752), .B1(n38057), .B2(n36659), .ZN(
        n7485) );
  OAI22_X1 U2130 ( .A1(n38060), .A2(n38759), .B1(n38057), .B2(n36661), .ZN(
        n7486) );
  OAI22_X1 U2131 ( .A1(n38060), .A2(n38766), .B1(n38057), .B2(n36663), .ZN(
        n7487) );
  OAI22_X1 U2132 ( .A1(n38060), .A2(n38773), .B1(n38057), .B2(n36665), .ZN(
        n7488) );
  OAI22_X1 U2133 ( .A1(n38060), .A2(n38780), .B1(n4668), .B2(n36667), .ZN(
        n7489) );
  OAI22_X1 U2134 ( .A1(n38061), .A2(n38787), .B1(n4668), .B2(n36669), .ZN(
        n7490) );
  OAI22_X1 U2135 ( .A1(n38061), .A2(n38794), .B1(n4668), .B2(n36671), .ZN(
        n7491) );
  OAI22_X1 U2136 ( .A1(n38061), .A2(n38801), .B1(n4668), .B2(n36673), .ZN(
        n7492) );
  OAI22_X1 U2137 ( .A1(n38061), .A2(n38808), .B1(n4668), .B2(n36675), .ZN(
        n7493) );
  OAI22_X1 U2138 ( .A1(n38061), .A2(n38815), .B1(n4668), .B2(n36677), .ZN(
        n7494) );
  OAI22_X1 U2139 ( .A1(n38062), .A2(n38822), .B1(n4668), .B2(n36679), .ZN(
        n7495) );
  OAI22_X1 U2140 ( .A1(n38062), .A2(n38829), .B1(n38057), .B2(n36681), .ZN(
        n7496) );
  OAI22_X1 U2141 ( .A1(n38062), .A2(n38836), .B1(n38057), .B2(n36683), .ZN(
        n7497) );
  OAI22_X1 U2142 ( .A1(n38062), .A2(n38843), .B1(n38057), .B2(n36685), .ZN(
        n7498) );
  OAI22_X1 U2143 ( .A1(n38079), .A2(n38681), .B1(n38078), .B2(n35929), .ZN(
        n7539) );
  OAI22_X1 U2144 ( .A1(n38079), .A2(n38688), .B1(n38078), .B2(n35933), .ZN(
        n7540) );
  OAI22_X1 U2145 ( .A1(n38079), .A2(n38695), .B1(n38078), .B2(n35937), .ZN(
        n7541) );
  OAI22_X1 U2146 ( .A1(n38079), .A2(n38702), .B1(n38078), .B2(n35941), .ZN(
        n7542) );
  OAI22_X1 U2147 ( .A1(n38079), .A2(n38709), .B1(n38078), .B2(n35945), .ZN(
        n7543) );
  OAI22_X1 U2148 ( .A1(n38080), .A2(n38716), .B1(n38078), .B2(n35949), .ZN(
        n7544) );
  OAI22_X1 U2149 ( .A1(n38080), .A2(n38723), .B1(n38078), .B2(n35953), .ZN(
        n7545) );
  OAI22_X1 U2150 ( .A1(n38080), .A2(n38730), .B1(n38078), .B2(n35957), .ZN(
        n7546) );
  OAI22_X1 U2151 ( .A1(n38080), .A2(n38737), .B1(n38078), .B2(n35961), .ZN(
        n7547) );
  OAI22_X1 U2152 ( .A1(n38080), .A2(n38744), .B1(n38078), .B2(n35965), .ZN(
        n7548) );
  OAI22_X1 U2153 ( .A1(n38081), .A2(n38751), .B1(n38078), .B2(n35969), .ZN(
        n7549) );
  OAI22_X1 U2154 ( .A1(n38081), .A2(n38758), .B1(n38078), .B2(n35973), .ZN(
        n7550) );
  OAI22_X1 U2155 ( .A1(n38081), .A2(n38765), .B1(n38078), .B2(n35977), .ZN(
        n7551) );
  OAI22_X1 U2156 ( .A1(n38081), .A2(n38772), .B1(n38078), .B2(n35981), .ZN(
        n7552) );
  OAI22_X1 U2157 ( .A1(n38081), .A2(n38779), .B1(n4598), .B2(n35985), .ZN(
        n7553) );
  OAI22_X1 U2158 ( .A1(n38082), .A2(n38786), .B1(n4598), .B2(n35989), .ZN(
        n7554) );
  OAI22_X1 U2159 ( .A1(n38082), .A2(n38793), .B1(n4598), .B2(n35993), .ZN(
        n7555) );
  OAI22_X1 U2160 ( .A1(n38082), .A2(n38800), .B1(n4598), .B2(n35997), .ZN(
        n7556) );
  OAI22_X1 U2161 ( .A1(n38082), .A2(n38807), .B1(n4598), .B2(n36001), .ZN(
        n7557) );
  OAI22_X1 U2162 ( .A1(n38082), .A2(n38814), .B1(n4598), .B2(n36005), .ZN(
        n7558) );
  OAI22_X1 U2163 ( .A1(n38083), .A2(n38821), .B1(n4598), .B2(n36009), .ZN(
        n7559) );
  OAI22_X1 U2164 ( .A1(n38083), .A2(n38828), .B1(n38078), .B2(n36013), .ZN(
        n7560) );
  OAI22_X1 U2165 ( .A1(n38083), .A2(n38835), .B1(n38078), .B2(n36017), .ZN(
        n7561) );
  OAI22_X1 U2166 ( .A1(n38083), .A2(n38842), .B1(n38078), .B2(n36021), .ZN(
        n7562) );
  OAI22_X1 U2167 ( .A1(n38091), .A2(n38681), .B1(n38090), .B2(n35519), .ZN(
        n7571) );
  OAI22_X1 U2168 ( .A1(n38091), .A2(n38688), .B1(n38090), .B2(n35521), .ZN(
        n7572) );
  OAI22_X1 U2169 ( .A1(n38091), .A2(n38695), .B1(n38090), .B2(n35523), .ZN(
        n7573) );
  OAI22_X1 U2170 ( .A1(n38091), .A2(n38702), .B1(n38090), .B2(n35525), .ZN(
        n7574) );
  OAI22_X1 U2171 ( .A1(n38091), .A2(n38709), .B1(n38090), .B2(n35527), .ZN(
        n7575) );
  OAI22_X1 U2172 ( .A1(n38092), .A2(n38716), .B1(n38090), .B2(n35529), .ZN(
        n7576) );
  OAI22_X1 U2173 ( .A1(n38092), .A2(n38723), .B1(n38090), .B2(n35531), .ZN(
        n7577) );
  OAI22_X1 U2174 ( .A1(n38092), .A2(n38730), .B1(n38090), .B2(n35533), .ZN(
        n7578) );
  OAI22_X1 U2175 ( .A1(n38092), .A2(n38737), .B1(n38090), .B2(n35535), .ZN(
        n7579) );
  OAI22_X1 U2176 ( .A1(n38092), .A2(n38744), .B1(n38090), .B2(n35537), .ZN(
        n7580) );
  OAI22_X1 U2177 ( .A1(n38093), .A2(n38751), .B1(n38090), .B2(n35539), .ZN(
        n7581) );
  OAI22_X1 U2178 ( .A1(n38093), .A2(n38758), .B1(n38090), .B2(n35541), .ZN(
        n7582) );
  OAI22_X1 U2179 ( .A1(n38093), .A2(n38765), .B1(n38090), .B2(n35543), .ZN(
        n7583) );
  OAI22_X1 U2180 ( .A1(n38093), .A2(n38772), .B1(n38090), .B2(n35545), .ZN(
        n7584) );
  OAI22_X1 U2181 ( .A1(n38093), .A2(n38779), .B1(n4563), .B2(n35547), .ZN(
        n7585) );
  OAI22_X1 U2182 ( .A1(n38094), .A2(n38786), .B1(n4563), .B2(n35549), .ZN(
        n7586) );
  OAI22_X1 U2183 ( .A1(n38094), .A2(n38793), .B1(n4563), .B2(n35551), .ZN(
        n7587) );
  OAI22_X1 U2184 ( .A1(n38094), .A2(n38800), .B1(n4563), .B2(n35553), .ZN(
        n7588) );
  OAI22_X1 U2185 ( .A1(n38094), .A2(n38807), .B1(n4563), .B2(n35555), .ZN(
        n7589) );
  OAI22_X1 U2186 ( .A1(n38094), .A2(n38814), .B1(n4563), .B2(n35557), .ZN(
        n7590) );
  OAI22_X1 U2187 ( .A1(n38095), .A2(n38821), .B1(n4563), .B2(n35559), .ZN(
        n7591) );
  OAI22_X1 U2188 ( .A1(n38095), .A2(n38828), .B1(n38090), .B2(n35561), .ZN(
        n7592) );
  OAI22_X1 U2189 ( .A1(n38095), .A2(n38835), .B1(n38090), .B2(n35563), .ZN(
        n7593) );
  OAI22_X1 U2190 ( .A1(n38095), .A2(n38842), .B1(n38090), .B2(n35565), .ZN(
        n7594) );
  OAI22_X1 U2191 ( .A1(n38112), .A2(n38681), .B1(n38111), .B2(n36270), .ZN(
        n7635) );
  OAI22_X1 U2192 ( .A1(n38112), .A2(n38688), .B1(n38111), .B2(n36271), .ZN(
        n7636) );
  OAI22_X1 U2193 ( .A1(n38112), .A2(n38695), .B1(n38111), .B2(n36272), .ZN(
        n7637) );
  OAI22_X1 U2194 ( .A1(n38112), .A2(n38702), .B1(n38111), .B2(n36273), .ZN(
        n7638) );
  OAI22_X1 U2195 ( .A1(n38112), .A2(n38709), .B1(n38111), .B2(n36274), .ZN(
        n7639) );
  OAI22_X1 U2196 ( .A1(n38113), .A2(n38716), .B1(n38111), .B2(n36275), .ZN(
        n7640) );
  OAI22_X1 U2197 ( .A1(n38113), .A2(n38723), .B1(n38111), .B2(n36276), .ZN(
        n7641) );
  OAI22_X1 U2198 ( .A1(n38113), .A2(n38730), .B1(n38111), .B2(n36277), .ZN(
        n7642) );
  OAI22_X1 U2199 ( .A1(n38113), .A2(n38737), .B1(n38111), .B2(n36278), .ZN(
        n7643) );
  OAI22_X1 U2200 ( .A1(n38113), .A2(n38744), .B1(n38111), .B2(n36279), .ZN(
        n7644) );
  OAI22_X1 U2201 ( .A1(n38114), .A2(n38751), .B1(n38111), .B2(n36280), .ZN(
        n7645) );
  OAI22_X1 U2202 ( .A1(n38114), .A2(n38758), .B1(n38111), .B2(n36281), .ZN(
        n7646) );
  OAI22_X1 U2203 ( .A1(n38114), .A2(n38765), .B1(n38111), .B2(n36282), .ZN(
        n7647) );
  OAI22_X1 U2204 ( .A1(n38114), .A2(n38772), .B1(n38111), .B2(n36283), .ZN(
        n7648) );
  OAI22_X1 U2205 ( .A1(n38114), .A2(n38779), .B1(n4493), .B2(n36284), .ZN(
        n7649) );
  OAI22_X1 U2206 ( .A1(n38115), .A2(n38786), .B1(n4493), .B2(n36285), .ZN(
        n7650) );
  OAI22_X1 U2207 ( .A1(n38115), .A2(n38793), .B1(n4493), .B2(n36286), .ZN(
        n7651) );
  OAI22_X1 U2208 ( .A1(n38115), .A2(n38800), .B1(n4493), .B2(n36287), .ZN(
        n7652) );
  OAI22_X1 U2209 ( .A1(n38115), .A2(n38807), .B1(n4493), .B2(n36288), .ZN(
        n7653) );
  OAI22_X1 U2210 ( .A1(n38115), .A2(n38814), .B1(n4493), .B2(n36289), .ZN(
        n7654) );
  OAI22_X1 U2211 ( .A1(n38116), .A2(n38821), .B1(n4493), .B2(n36290), .ZN(
        n7655) );
  OAI22_X1 U2212 ( .A1(n38116), .A2(n38828), .B1(n38111), .B2(n36291), .ZN(
        n7656) );
  OAI22_X1 U2213 ( .A1(n38116), .A2(n38835), .B1(n38111), .B2(n36292), .ZN(
        n7657) );
  OAI22_X1 U2214 ( .A1(n38116), .A2(n38842), .B1(n38111), .B2(n36293), .ZN(
        n7658) );
  OAI22_X1 U2215 ( .A1(n38133), .A2(n38681), .B1(n38132), .B2(n35758), .ZN(
        n7699) );
  OAI22_X1 U2216 ( .A1(n38133), .A2(n38688), .B1(n38132), .B2(n35759), .ZN(
        n7700) );
  OAI22_X1 U2217 ( .A1(n38133), .A2(n38695), .B1(n38132), .B2(n35760), .ZN(
        n7701) );
  OAI22_X1 U2218 ( .A1(n38133), .A2(n38702), .B1(n38132), .B2(n35761), .ZN(
        n7702) );
  OAI22_X1 U2219 ( .A1(n38133), .A2(n38709), .B1(n38132), .B2(n35762), .ZN(
        n7703) );
  OAI22_X1 U2220 ( .A1(n38134), .A2(n38716), .B1(n38132), .B2(n35763), .ZN(
        n7704) );
  OAI22_X1 U2221 ( .A1(n38134), .A2(n38723), .B1(n38132), .B2(n35764), .ZN(
        n7705) );
  OAI22_X1 U2222 ( .A1(n38134), .A2(n38730), .B1(n38132), .B2(n35765), .ZN(
        n7706) );
  OAI22_X1 U2223 ( .A1(n38134), .A2(n38737), .B1(n38132), .B2(n35766), .ZN(
        n7707) );
  OAI22_X1 U2224 ( .A1(n38134), .A2(n38744), .B1(n38132), .B2(n35767), .ZN(
        n7708) );
  OAI22_X1 U2225 ( .A1(n38135), .A2(n38751), .B1(n38132), .B2(n35768), .ZN(
        n7709) );
  OAI22_X1 U2226 ( .A1(n38135), .A2(n38758), .B1(n38132), .B2(n35769), .ZN(
        n7710) );
  OAI22_X1 U2227 ( .A1(n38135), .A2(n38765), .B1(n38132), .B2(n35770), .ZN(
        n7711) );
  OAI22_X1 U2228 ( .A1(n38135), .A2(n38772), .B1(n38132), .B2(n35771), .ZN(
        n7712) );
  OAI22_X1 U2229 ( .A1(n38135), .A2(n38779), .B1(n4423), .B2(n35772), .ZN(
        n7713) );
  OAI22_X1 U2230 ( .A1(n38136), .A2(n38786), .B1(n4423), .B2(n35773), .ZN(
        n7714) );
  OAI22_X1 U2231 ( .A1(n38136), .A2(n38793), .B1(n4423), .B2(n35774), .ZN(
        n7715) );
  OAI22_X1 U2232 ( .A1(n38136), .A2(n38800), .B1(n4423), .B2(n35775), .ZN(
        n7716) );
  OAI22_X1 U2233 ( .A1(n38136), .A2(n38807), .B1(n4423), .B2(n35776), .ZN(
        n7717) );
  OAI22_X1 U2234 ( .A1(n38136), .A2(n38814), .B1(n4423), .B2(n35777), .ZN(
        n7718) );
  OAI22_X1 U2235 ( .A1(n38137), .A2(n38821), .B1(n4423), .B2(n35778), .ZN(
        n7719) );
  OAI22_X1 U2236 ( .A1(n38137), .A2(n38828), .B1(n38132), .B2(n35779), .ZN(
        n7720) );
  OAI22_X1 U2237 ( .A1(n38137), .A2(n38835), .B1(n38132), .B2(n35780), .ZN(
        n7721) );
  OAI22_X1 U2238 ( .A1(n38137), .A2(n38842), .B1(n38132), .B2(n35781), .ZN(
        n7722) );
  OAI22_X1 U2239 ( .A1(n38145), .A2(n38681), .B1(n38144), .B2(n36590), .ZN(
        n7731) );
  OAI22_X1 U2240 ( .A1(n38145), .A2(n38688), .B1(n38144), .B2(n36592), .ZN(
        n7732) );
  OAI22_X1 U2241 ( .A1(n38145), .A2(n38695), .B1(n38144), .B2(n36594), .ZN(
        n7733) );
  OAI22_X1 U2242 ( .A1(n38145), .A2(n38702), .B1(n38144), .B2(n36596), .ZN(
        n7734) );
  OAI22_X1 U2243 ( .A1(n38145), .A2(n38709), .B1(n38144), .B2(n36598), .ZN(
        n7735) );
  OAI22_X1 U2244 ( .A1(n38146), .A2(n38716), .B1(n38144), .B2(n36600), .ZN(
        n7736) );
  OAI22_X1 U2245 ( .A1(n38146), .A2(n38723), .B1(n38144), .B2(n36602), .ZN(
        n7737) );
  OAI22_X1 U2246 ( .A1(n38146), .A2(n38730), .B1(n38144), .B2(n36604), .ZN(
        n7738) );
  OAI22_X1 U2247 ( .A1(n38146), .A2(n38737), .B1(n38144), .B2(n36606), .ZN(
        n7739) );
  OAI22_X1 U2248 ( .A1(n38146), .A2(n38744), .B1(n38144), .B2(n36608), .ZN(
        n7740) );
  OAI22_X1 U2249 ( .A1(n38147), .A2(n38751), .B1(n38144), .B2(n36610), .ZN(
        n7741) );
  OAI22_X1 U2250 ( .A1(n38147), .A2(n38758), .B1(n38144), .B2(n36612), .ZN(
        n7742) );
  OAI22_X1 U2251 ( .A1(n38147), .A2(n38765), .B1(n38144), .B2(n36614), .ZN(
        n7743) );
  OAI22_X1 U2252 ( .A1(n38147), .A2(n38772), .B1(n38144), .B2(n36616), .ZN(
        n7744) );
  OAI22_X1 U2253 ( .A1(n38147), .A2(n38779), .B1(n4388), .B2(n36618), .ZN(
        n7745) );
  OAI22_X1 U2254 ( .A1(n38148), .A2(n38786), .B1(n4388), .B2(n36620), .ZN(
        n7746) );
  OAI22_X1 U2255 ( .A1(n38148), .A2(n38793), .B1(n4388), .B2(n36622), .ZN(
        n7747) );
  OAI22_X1 U2256 ( .A1(n38148), .A2(n38800), .B1(n4388), .B2(n36624), .ZN(
        n7748) );
  OAI22_X1 U2257 ( .A1(n38148), .A2(n38807), .B1(n4388), .B2(n36626), .ZN(
        n7749) );
  OAI22_X1 U2258 ( .A1(n38148), .A2(n38814), .B1(n4388), .B2(n36628), .ZN(
        n7750) );
  OAI22_X1 U2259 ( .A1(n38149), .A2(n38821), .B1(n4388), .B2(n36630), .ZN(
        n7751) );
  OAI22_X1 U2260 ( .A1(n38149), .A2(n38828), .B1(n38144), .B2(n36632), .ZN(
        n7752) );
  OAI22_X1 U2261 ( .A1(n38149), .A2(n38835), .B1(n38144), .B2(n36634), .ZN(
        n7753) );
  OAI22_X1 U2262 ( .A1(n38149), .A2(n38842), .B1(n38144), .B2(n36636), .ZN(
        n7754) );
  OAI22_X1 U2263 ( .A1(n38166), .A2(n38681), .B1(n38165), .B2(n36126), .ZN(
        n7795) );
  OAI22_X1 U2264 ( .A1(n38166), .A2(n38688), .B1(n38165), .B2(n36128), .ZN(
        n7796) );
  OAI22_X1 U2265 ( .A1(n38166), .A2(n38695), .B1(n38165), .B2(n36130), .ZN(
        n7797) );
  OAI22_X1 U2266 ( .A1(n38166), .A2(n38702), .B1(n38165), .B2(n36132), .ZN(
        n7798) );
  OAI22_X1 U2267 ( .A1(n38166), .A2(n38709), .B1(n38165), .B2(n36134), .ZN(
        n7799) );
  OAI22_X1 U2268 ( .A1(n38167), .A2(n38716), .B1(n38165), .B2(n36136), .ZN(
        n7800) );
  OAI22_X1 U2269 ( .A1(n38167), .A2(n38723), .B1(n38165), .B2(n36138), .ZN(
        n7801) );
  OAI22_X1 U2270 ( .A1(n38167), .A2(n38730), .B1(n38165), .B2(n36140), .ZN(
        n7802) );
  OAI22_X1 U2271 ( .A1(n38167), .A2(n38737), .B1(n38165), .B2(n36142), .ZN(
        n7803) );
  OAI22_X1 U2272 ( .A1(n38167), .A2(n38744), .B1(n38165), .B2(n36144), .ZN(
        n7804) );
  OAI22_X1 U2273 ( .A1(n38168), .A2(n38751), .B1(n38165), .B2(n36146), .ZN(
        n7805) );
  OAI22_X1 U2274 ( .A1(n38168), .A2(n38758), .B1(n38165), .B2(n36148), .ZN(
        n7806) );
  OAI22_X1 U2275 ( .A1(n38168), .A2(n38765), .B1(n38165), .B2(n36150), .ZN(
        n7807) );
  OAI22_X1 U2276 ( .A1(n38168), .A2(n38772), .B1(n38165), .B2(n36152), .ZN(
        n7808) );
  OAI22_X1 U2277 ( .A1(n38168), .A2(n38779), .B1(n4318), .B2(n36154), .ZN(
        n7809) );
  OAI22_X1 U2278 ( .A1(n38169), .A2(n38786), .B1(n4318), .B2(n36156), .ZN(
        n7810) );
  OAI22_X1 U2279 ( .A1(n38169), .A2(n38793), .B1(n4318), .B2(n36158), .ZN(
        n7811) );
  OAI22_X1 U2280 ( .A1(n38169), .A2(n38800), .B1(n4318), .B2(n36160), .ZN(
        n7812) );
  OAI22_X1 U2281 ( .A1(n38169), .A2(n38807), .B1(n4318), .B2(n36162), .ZN(
        n7813) );
  OAI22_X1 U2282 ( .A1(n38169), .A2(n38814), .B1(n4318), .B2(n36164), .ZN(
        n7814) );
  OAI22_X1 U2283 ( .A1(n38170), .A2(n38821), .B1(n4318), .B2(n36166), .ZN(
        n7815) );
  OAI22_X1 U2284 ( .A1(n38170), .A2(n38828), .B1(n38165), .B2(n36168), .ZN(
        n7816) );
  OAI22_X1 U2285 ( .A1(n38170), .A2(n38835), .B1(n38165), .B2(n36170), .ZN(
        n7817) );
  OAI22_X1 U2286 ( .A1(n38170), .A2(n38842), .B1(n38165), .B2(n36172), .ZN(
        n7818) );
  OAI22_X1 U2287 ( .A1(n38178), .A2(n38681), .B1(n38177), .B2(n35416), .ZN(
        n7827) );
  OAI22_X1 U2288 ( .A1(n38178), .A2(n38688), .B1(n38177), .B2(n35420), .ZN(
        n7828) );
  OAI22_X1 U2289 ( .A1(n38178), .A2(n38695), .B1(n38177), .B2(n35424), .ZN(
        n7829) );
  OAI22_X1 U2290 ( .A1(n38178), .A2(n38702), .B1(n38177), .B2(n35428), .ZN(
        n7830) );
  OAI22_X1 U2291 ( .A1(n38178), .A2(n38709), .B1(n38177), .B2(n35432), .ZN(
        n7831) );
  OAI22_X1 U2292 ( .A1(n38179), .A2(n38716), .B1(n38177), .B2(n35436), .ZN(
        n7832) );
  OAI22_X1 U2293 ( .A1(n38179), .A2(n38723), .B1(n38177), .B2(n35440), .ZN(
        n7833) );
  OAI22_X1 U2294 ( .A1(n38179), .A2(n38730), .B1(n38177), .B2(n35444), .ZN(
        n7834) );
  OAI22_X1 U2295 ( .A1(n38179), .A2(n38737), .B1(n38177), .B2(n35448), .ZN(
        n7835) );
  OAI22_X1 U2296 ( .A1(n38179), .A2(n38744), .B1(n38177), .B2(n35452), .ZN(
        n7836) );
  OAI22_X1 U2297 ( .A1(n38180), .A2(n38751), .B1(n38177), .B2(n35456), .ZN(
        n7837) );
  OAI22_X1 U2298 ( .A1(n38180), .A2(n38758), .B1(n38177), .B2(n35460), .ZN(
        n7838) );
  OAI22_X1 U2299 ( .A1(n38180), .A2(n38765), .B1(n38177), .B2(n35464), .ZN(
        n7839) );
  OAI22_X1 U2300 ( .A1(n38180), .A2(n38772), .B1(n38177), .B2(n35468), .ZN(
        n7840) );
  OAI22_X1 U2301 ( .A1(n38180), .A2(n38779), .B1(n4283), .B2(n35472), .ZN(
        n7841) );
  OAI22_X1 U2302 ( .A1(n38181), .A2(n38786), .B1(n4283), .B2(n35476), .ZN(
        n7842) );
  OAI22_X1 U2303 ( .A1(n38181), .A2(n38793), .B1(n4283), .B2(n35480), .ZN(
        n7843) );
  OAI22_X1 U2304 ( .A1(n38181), .A2(n38800), .B1(n4283), .B2(n35484), .ZN(
        n7844) );
  OAI22_X1 U2305 ( .A1(n38181), .A2(n38807), .B1(n4283), .B2(n35488), .ZN(
        n7845) );
  OAI22_X1 U2306 ( .A1(n38181), .A2(n38814), .B1(n4283), .B2(n35492), .ZN(
        n7846) );
  OAI22_X1 U2307 ( .A1(n38182), .A2(n38821), .B1(n4283), .B2(n35496), .ZN(
        n7847) );
  OAI22_X1 U2308 ( .A1(n38182), .A2(n38828), .B1(n38177), .B2(n35500), .ZN(
        n7848) );
  OAI22_X1 U2309 ( .A1(n38182), .A2(n38835), .B1(n38177), .B2(n35504), .ZN(
        n7849) );
  OAI22_X1 U2310 ( .A1(n38182), .A2(n38842), .B1(n38177), .B2(n35508), .ZN(
        n7850) );
  OAI22_X1 U2311 ( .A1(n38199), .A2(n38680), .B1(n38198), .B2(n36542), .ZN(
        n7891) );
  OAI22_X1 U2312 ( .A1(n38199), .A2(n38687), .B1(n38198), .B2(n36544), .ZN(
        n7892) );
  OAI22_X1 U2313 ( .A1(n38199), .A2(n38694), .B1(n38198), .B2(n36546), .ZN(
        n7893) );
  OAI22_X1 U2314 ( .A1(n38199), .A2(n38701), .B1(n38198), .B2(n36548), .ZN(
        n7894) );
  OAI22_X1 U2315 ( .A1(n38199), .A2(n38708), .B1(n38198), .B2(n36550), .ZN(
        n7895) );
  OAI22_X1 U2316 ( .A1(n38200), .A2(n38715), .B1(n38198), .B2(n36552), .ZN(
        n7896) );
  OAI22_X1 U2317 ( .A1(n38200), .A2(n38722), .B1(n38198), .B2(n36554), .ZN(
        n7897) );
  OAI22_X1 U2318 ( .A1(n38200), .A2(n38729), .B1(n38198), .B2(n36556), .ZN(
        n7898) );
  OAI22_X1 U2319 ( .A1(n38200), .A2(n38736), .B1(n38198), .B2(n36558), .ZN(
        n7899) );
  OAI22_X1 U2320 ( .A1(n38200), .A2(n38743), .B1(n38198), .B2(n36560), .ZN(
        n7900) );
  OAI22_X1 U2321 ( .A1(n38201), .A2(n38750), .B1(n38198), .B2(n36562), .ZN(
        n7901) );
  OAI22_X1 U2322 ( .A1(n38201), .A2(n38757), .B1(n38198), .B2(n36564), .ZN(
        n7902) );
  OAI22_X1 U2323 ( .A1(n38201), .A2(n38764), .B1(n38198), .B2(n36566), .ZN(
        n7903) );
  OAI22_X1 U2324 ( .A1(n38201), .A2(n38771), .B1(n38198), .B2(n36568), .ZN(
        n7904) );
  OAI22_X1 U2325 ( .A1(n38201), .A2(n38778), .B1(n4213), .B2(n36570), .ZN(
        n7905) );
  OAI22_X1 U2326 ( .A1(n38202), .A2(n38785), .B1(n4213), .B2(n36572), .ZN(
        n7906) );
  OAI22_X1 U2327 ( .A1(n38202), .A2(n38792), .B1(n4213), .B2(n36574), .ZN(
        n7907) );
  OAI22_X1 U2328 ( .A1(n38202), .A2(n38799), .B1(n4213), .B2(n36576), .ZN(
        n7908) );
  OAI22_X1 U2329 ( .A1(n38202), .A2(n38806), .B1(n4213), .B2(n36578), .ZN(
        n7909) );
  OAI22_X1 U2330 ( .A1(n38202), .A2(n38813), .B1(n4213), .B2(n36580), .ZN(
        n7910) );
  OAI22_X1 U2331 ( .A1(n38203), .A2(n38820), .B1(n4213), .B2(n36582), .ZN(
        n7911) );
  OAI22_X1 U2332 ( .A1(n38203), .A2(n38827), .B1(n38198), .B2(n36584), .ZN(
        n7912) );
  OAI22_X1 U2333 ( .A1(n38203), .A2(n38834), .B1(n38198), .B2(n36586), .ZN(
        n7913) );
  OAI22_X1 U2334 ( .A1(n38203), .A2(n38841), .B1(n38198), .B2(n36588), .ZN(
        n7914) );
  OAI22_X1 U2335 ( .A1(n38220), .A2(n38680), .B1(n38219), .B2(n36079), .ZN(
        n7955) );
  OAI22_X1 U2336 ( .A1(n38220), .A2(n38687), .B1(n38219), .B2(n36081), .ZN(
        n7956) );
  OAI22_X1 U2337 ( .A1(n38220), .A2(n38694), .B1(n38219), .B2(n36083), .ZN(
        n7957) );
  OAI22_X1 U2338 ( .A1(n38220), .A2(n38701), .B1(n38219), .B2(n36085), .ZN(
        n7958) );
  OAI22_X1 U2339 ( .A1(n38220), .A2(n38708), .B1(n38219), .B2(n36087), .ZN(
        n7959) );
  OAI22_X1 U2340 ( .A1(n38221), .A2(n38715), .B1(n38219), .B2(n36089), .ZN(
        n7960) );
  OAI22_X1 U2341 ( .A1(n38221), .A2(n38722), .B1(n38219), .B2(n36091), .ZN(
        n7961) );
  OAI22_X1 U2342 ( .A1(n38221), .A2(n38729), .B1(n38219), .B2(n36093), .ZN(
        n7962) );
  OAI22_X1 U2343 ( .A1(n38221), .A2(n38736), .B1(n38219), .B2(n36095), .ZN(
        n7963) );
  OAI22_X1 U2344 ( .A1(n38221), .A2(n38743), .B1(n38219), .B2(n36097), .ZN(
        n7964) );
  OAI22_X1 U2345 ( .A1(n38222), .A2(n38750), .B1(n38219), .B2(n36099), .ZN(
        n7965) );
  OAI22_X1 U2346 ( .A1(n38222), .A2(n38757), .B1(n38219), .B2(n36101), .ZN(
        n7966) );
  OAI22_X1 U2347 ( .A1(n38222), .A2(n38764), .B1(n38219), .B2(n36103), .ZN(
        n7967) );
  OAI22_X1 U2348 ( .A1(n38222), .A2(n38771), .B1(n38219), .B2(n36105), .ZN(
        n7968) );
  OAI22_X1 U2349 ( .A1(n38222), .A2(n38778), .B1(n4140), .B2(n36107), .ZN(
        n7969) );
  OAI22_X1 U2350 ( .A1(n38223), .A2(n38785), .B1(n4140), .B2(n36109), .ZN(
        n7970) );
  OAI22_X1 U2351 ( .A1(n38223), .A2(n38792), .B1(n4140), .B2(n36111), .ZN(
        n7971) );
  OAI22_X1 U2352 ( .A1(n38223), .A2(n38799), .B1(n4140), .B2(n36113), .ZN(
        n7972) );
  OAI22_X1 U2353 ( .A1(n38223), .A2(n38806), .B1(n4140), .B2(n36115), .ZN(
        n7973) );
  OAI22_X1 U2354 ( .A1(n38223), .A2(n38813), .B1(n4140), .B2(n36117), .ZN(
        n7974) );
  OAI22_X1 U2355 ( .A1(n38224), .A2(n38820), .B1(n4140), .B2(n36119), .ZN(
        n7975) );
  OAI22_X1 U2356 ( .A1(n38224), .A2(n38827), .B1(n38219), .B2(n36121), .ZN(
        n7976) );
  OAI22_X1 U2357 ( .A1(n38224), .A2(n38834), .B1(n38219), .B2(n36123), .ZN(
        n7977) );
  OAI22_X1 U2358 ( .A1(n38224), .A2(n38841), .B1(n38219), .B2(n36125), .ZN(
        n7978) );
  OAI22_X1 U2359 ( .A1(n38232), .A2(n38680), .B1(n38231), .B2(n35615), .ZN(
        n7987) );
  OAI22_X1 U2360 ( .A1(n38232), .A2(n38687), .B1(n38231), .B2(n35617), .ZN(
        n7988) );
  OAI22_X1 U2361 ( .A1(n38232), .A2(n38694), .B1(n38231), .B2(n35619), .ZN(
        n7989) );
  OAI22_X1 U2362 ( .A1(n38232), .A2(n38701), .B1(n38231), .B2(n35621), .ZN(
        n7990) );
  OAI22_X1 U2363 ( .A1(n38232), .A2(n38708), .B1(n38231), .B2(n35623), .ZN(
        n7991) );
  OAI22_X1 U2364 ( .A1(n38233), .A2(n38715), .B1(n38231), .B2(n35625), .ZN(
        n7992) );
  OAI22_X1 U2365 ( .A1(n38233), .A2(n38722), .B1(n38231), .B2(n35627), .ZN(
        n7993) );
  OAI22_X1 U2366 ( .A1(n38233), .A2(n38729), .B1(n38231), .B2(n35629), .ZN(
        n7994) );
  OAI22_X1 U2367 ( .A1(n38233), .A2(n38736), .B1(n38231), .B2(n35631), .ZN(
        n7995) );
  OAI22_X1 U2368 ( .A1(n38233), .A2(n38743), .B1(n38231), .B2(n35633), .ZN(
        n7996) );
  OAI22_X1 U2369 ( .A1(n38234), .A2(n38750), .B1(n38231), .B2(n35635), .ZN(
        n7997) );
  OAI22_X1 U2370 ( .A1(n38234), .A2(n38757), .B1(n38231), .B2(n35637), .ZN(
        n7998) );
  OAI22_X1 U2371 ( .A1(n38234), .A2(n38764), .B1(n38231), .B2(n35639), .ZN(
        n7999) );
  OAI22_X1 U2372 ( .A1(n38234), .A2(n38771), .B1(n38231), .B2(n35641), .ZN(
        n8000) );
  OAI22_X1 U2373 ( .A1(n38234), .A2(n38778), .B1(n4076), .B2(n35643), .ZN(
        n8001) );
  OAI22_X1 U2374 ( .A1(n38235), .A2(n38785), .B1(n4076), .B2(n35645), .ZN(
        n8002) );
  OAI22_X1 U2375 ( .A1(n38235), .A2(n38792), .B1(n4076), .B2(n35647), .ZN(
        n8003) );
  OAI22_X1 U2376 ( .A1(n38235), .A2(n38799), .B1(n4076), .B2(n35649), .ZN(
        n8004) );
  OAI22_X1 U2377 ( .A1(n38235), .A2(n38806), .B1(n4076), .B2(n35651), .ZN(
        n8005) );
  OAI22_X1 U2378 ( .A1(n38235), .A2(n38813), .B1(n4076), .B2(n35653), .ZN(
        n8006) );
  OAI22_X1 U2379 ( .A1(n38236), .A2(n38820), .B1(n4076), .B2(n35655), .ZN(
        n8007) );
  OAI22_X1 U2380 ( .A1(n38236), .A2(n38827), .B1(n38231), .B2(n35657), .ZN(
        n8008) );
  OAI22_X1 U2381 ( .A1(n38236), .A2(n38834), .B1(n38231), .B2(n35659), .ZN(
        n8009) );
  OAI22_X1 U2382 ( .A1(n38236), .A2(n38841), .B1(n38231), .B2(n35661), .ZN(
        n8010) );
  OAI22_X1 U2383 ( .A1(n38253), .A2(n38680), .B1(n38252), .B2(n36441), .ZN(
        n8051) );
  OAI22_X1 U2384 ( .A1(n38253), .A2(n38687), .B1(n38252), .B2(n36445), .ZN(
        n8052) );
  OAI22_X1 U2385 ( .A1(n38253), .A2(n38694), .B1(n38252), .B2(n36449), .ZN(
        n8053) );
  OAI22_X1 U2386 ( .A1(n38253), .A2(n38701), .B1(n38252), .B2(n36453), .ZN(
        n8054) );
  OAI22_X1 U2387 ( .A1(n38253), .A2(n38708), .B1(n38252), .B2(n36457), .ZN(
        n8055) );
  OAI22_X1 U2388 ( .A1(n38254), .A2(n38715), .B1(n38252), .B2(n36461), .ZN(
        n8056) );
  OAI22_X1 U2389 ( .A1(n38254), .A2(n38722), .B1(n38252), .B2(n36465), .ZN(
        n8057) );
  OAI22_X1 U2390 ( .A1(n38254), .A2(n38729), .B1(n38252), .B2(n36469), .ZN(
        n8058) );
  OAI22_X1 U2391 ( .A1(n38254), .A2(n38736), .B1(n38252), .B2(n36473), .ZN(
        n8059) );
  OAI22_X1 U2392 ( .A1(n38254), .A2(n38743), .B1(n38252), .B2(n36477), .ZN(
        n8060) );
  OAI22_X1 U2393 ( .A1(n38255), .A2(n38750), .B1(n38252), .B2(n36481), .ZN(
        n8061) );
  OAI22_X1 U2394 ( .A1(n38255), .A2(n38757), .B1(n38252), .B2(n36485), .ZN(
        n8062) );
  OAI22_X1 U2395 ( .A1(n38255), .A2(n38764), .B1(n38252), .B2(n36489), .ZN(
        n8063) );
  OAI22_X1 U2396 ( .A1(n38255), .A2(n38771), .B1(n38252), .B2(n36493), .ZN(
        n8064) );
  OAI22_X1 U2397 ( .A1(n38255), .A2(n38778), .B1(n4006), .B2(n36497), .ZN(
        n8065) );
  OAI22_X1 U2398 ( .A1(n38256), .A2(n38785), .B1(n4006), .B2(n36501), .ZN(
        n8066) );
  OAI22_X1 U2399 ( .A1(n38256), .A2(n38792), .B1(n4006), .B2(n36505), .ZN(
        n8067) );
  OAI22_X1 U2400 ( .A1(n38256), .A2(n38799), .B1(n4006), .B2(n36509), .ZN(
        n8068) );
  OAI22_X1 U2401 ( .A1(n38256), .A2(n38806), .B1(n4006), .B2(n36513), .ZN(
        n8069) );
  OAI22_X1 U2402 ( .A1(n38256), .A2(n38813), .B1(n4006), .B2(n36517), .ZN(
        n8070) );
  OAI22_X1 U2403 ( .A1(n38257), .A2(n38820), .B1(n4006), .B2(n36521), .ZN(
        n8071) );
  OAI22_X1 U2404 ( .A1(n38257), .A2(n38827), .B1(n38252), .B2(n36525), .ZN(
        n8072) );
  OAI22_X1 U2405 ( .A1(n38257), .A2(n38834), .B1(n38252), .B2(n36529), .ZN(
        n8073) );
  OAI22_X1 U2406 ( .A1(n38257), .A2(n38841), .B1(n38252), .B2(n36533), .ZN(
        n8074) );
  OAI22_X1 U2407 ( .A1(n38274), .A2(n38680), .B1(n38273), .B2(n36031), .ZN(
        n8115) );
  OAI22_X1 U2408 ( .A1(n38274), .A2(n38687), .B1(n38273), .B2(n36033), .ZN(
        n8116) );
  OAI22_X1 U2409 ( .A1(n38274), .A2(n38694), .B1(n38273), .B2(n36035), .ZN(
        n8117) );
  OAI22_X1 U2410 ( .A1(n38274), .A2(n38701), .B1(n38273), .B2(n36037), .ZN(
        n8118) );
  OAI22_X1 U2411 ( .A1(n38274), .A2(n38708), .B1(n38273), .B2(n36039), .ZN(
        n8119) );
  OAI22_X1 U2412 ( .A1(n38275), .A2(n38715), .B1(n38273), .B2(n36041), .ZN(
        n8120) );
  OAI22_X1 U2413 ( .A1(n38275), .A2(n38722), .B1(n38273), .B2(n36043), .ZN(
        n8121) );
  OAI22_X1 U2414 ( .A1(n38275), .A2(n38729), .B1(n38273), .B2(n36045), .ZN(
        n8122) );
  OAI22_X1 U2415 ( .A1(n38275), .A2(n38736), .B1(n38273), .B2(n36047), .ZN(
        n8123) );
  OAI22_X1 U2416 ( .A1(n38275), .A2(n38743), .B1(n38273), .B2(n36049), .ZN(
        n8124) );
  OAI22_X1 U2417 ( .A1(n38276), .A2(n38750), .B1(n38273), .B2(n36051), .ZN(
        n8125) );
  OAI22_X1 U2418 ( .A1(n38276), .A2(n38757), .B1(n38273), .B2(n36053), .ZN(
        n8126) );
  OAI22_X1 U2419 ( .A1(n38276), .A2(n38764), .B1(n38273), .B2(n36055), .ZN(
        n8127) );
  OAI22_X1 U2420 ( .A1(n38276), .A2(n38771), .B1(n38273), .B2(n36057), .ZN(
        n8128) );
  OAI22_X1 U2421 ( .A1(n38276), .A2(n38778), .B1(n3936), .B2(n36059), .ZN(
        n8129) );
  OAI22_X1 U2422 ( .A1(n38277), .A2(n38785), .B1(n3936), .B2(n36061), .ZN(
        n8130) );
  OAI22_X1 U2423 ( .A1(n38277), .A2(n38792), .B1(n3936), .B2(n36063), .ZN(
        n8131) );
  OAI22_X1 U2424 ( .A1(n38277), .A2(n38799), .B1(n3936), .B2(n36065), .ZN(
        n8132) );
  OAI22_X1 U2425 ( .A1(n38277), .A2(n38806), .B1(n3936), .B2(n36067), .ZN(
        n8133) );
  OAI22_X1 U2426 ( .A1(n38277), .A2(n38813), .B1(n3936), .B2(n36069), .ZN(
        n8134) );
  OAI22_X1 U2427 ( .A1(n38278), .A2(n38820), .B1(n3936), .B2(n36071), .ZN(
        n8135) );
  OAI22_X1 U2428 ( .A1(n38278), .A2(n38827), .B1(n38273), .B2(n36073), .ZN(
        n8136) );
  OAI22_X1 U2429 ( .A1(n38278), .A2(n38834), .B1(n38273), .B2(n36075), .ZN(
        n8137) );
  OAI22_X1 U2430 ( .A1(n38278), .A2(n38841), .B1(n38273), .B2(n36077), .ZN(
        n8138) );
  OAI22_X1 U2431 ( .A1(n38286), .A2(n38680), .B1(n38285), .B2(n35246), .ZN(
        n8147) );
  OAI22_X1 U2432 ( .A1(n38286), .A2(n38687), .B1(n38285), .B2(n35247), .ZN(
        n8148) );
  OAI22_X1 U2433 ( .A1(n38286), .A2(n38694), .B1(n38285), .B2(n35248), .ZN(
        n8149) );
  OAI22_X1 U2434 ( .A1(n38286), .A2(n38701), .B1(n38285), .B2(n35249), .ZN(
        n8150) );
  OAI22_X1 U2435 ( .A1(n38286), .A2(n38708), .B1(n38285), .B2(n35250), .ZN(
        n8151) );
  OAI22_X1 U2436 ( .A1(n38287), .A2(n38715), .B1(n38285), .B2(n35251), .ZN(
        n8152) );
  OAI22_X1 U2437 ( .A1(n38287), .A2(n38722), .B1(n38285), .B2(n35252), .ZN(
        n8153) );
  OAI22_X1 U2438 ( .A1(n38287), .A2(n38729), .B1(n38285), .B2(n35253), .ZN(
        n8154) );
  OAI22_X1 U2439 ( .A1(n38287), .A2(n38736), .B1(n38285), .B2(n35254), .ZN(
        n8155) );
  OAI22_X1 U2440 ( .A1(n38287), .A2(n38743), .B1(n38285), .B2(n35255), .ZN(
        n8156) );
  OAI22_X1 U2441 ( .A1(n38288), .A2(n38750), .B1(n38285), .B2(n35256), .ZN(
        n8157) );
  OAI22_X1 U2442 ( .A1(n38288), .A2(n38757), .B1(n38285), .B2(n35257), .ZN(
        n8158) );
  OAI22_X1 U2443 ( .A1(n38288), .A2(n38764), .B1(n38285), .B2(n35258), .ZN(
        n8159) );
  OAI22_X1 U2444 ( .A1(n38288), .A2(n38771), .B1(n38285), .B2(n35259), .ZN(
        n8160) );
  OAI22_X1 U2445 ( .A1(n38288), .A2(n38778), .B1(n3901), .B2(n35260), .ZN(
        n8161) );
  OAI22_X1 U2446 ( .A1(n38289), .A2(n38785), .B1(n3901), .B2(n35261), .ZN(
        n8162) );
  OAI22_X1 U2447 ( .A1(n38289), .A2(n38792), .B1(n3901), .B2(n35262), .ZN(
        n8163) );
  OAI22_X1 U2448 ( .A1(n38289), .A2(n38799), .B1(n3901), .B2(n35263), .ZN(
        n8164) );
  OAI22_X1 U2449 ( .A1(n38289), .A2(n38806), .B1(n3901), .B2(n35264), .ZN(
        n8165) );
  OAI22_X1 U2450 ( .A1(n38289), .A2(n38813), .B1(n3901), .B2(n35265), .ZN(
        n8166) );
  OAI22_X1 U2451 ( .A1(n38290), .A2(n38820), .B1(n3901), .B2(n35266), .ZN(
        n8167) );
  OAI22_X1 U2452 ( .A1(n38290), .A2(n38827), .B1(n38285), .B2(n35267), .ZN(
        n8168) );
  OAI22_X1 U2453 ( .A1(n38290), .A2(n38834), .B1(n38285), .B2(n35268), .ZN(
        n8169) );
  OAI22_X1 U2454 ( .A1(n38290), .A2(n38841), .B1(n38285), .B2(n35269), .ZN(
        n8170) );
  OAI22_X1 U2455 ( .A1(n38307), .A2(n38680), .B1(n38306), .B2(n36294), .ZN(
        n8211) );
  OAI22_X1 U2456 ( .A1(n38307), .A2(n38687), .B1(n38306), .B2(n36295), .ZN(
        n8212) );
  OAI22_X1 U2457 ( .A1(n38307), .A2(n38694), .B1(n38306), .B2(n36296), .ZN(
        n8213) );
  OAI22_X1 U2458 ( .A1(n38307), .A2(n38701), .B1(n38306), .B2(n36297), .ZN(
        n8214) );
  OAI22_X1 U2459 ( .A1(n38307), .A2(n38708), .B1(n38306), .B2(n36298), .ZN(
        n8215) );
  OAI22_X1 U2460 ( .A1(n38308), .A2(n38715), .B1(n38306), .B2(n36299), .ZN(
        n8216) );
  OAI22_X1 U2461 ( .A1(n38308), .A2(n38722), .B1(n38306), .B2(n36300), .ZN(
        n8217) );
  OAI22_X1 U2462 ( .A1(n38308), .A2(n38729), .B1(n38306), .B2(n36301), .ZN(
        n8218) );
  OAI22_X1 U2463 ( .A1(n38308), .A2(n38736), .B1(n38306), .B2(n36302), .ZN(
        n8219) );
  OAI22_X1 U2464 ( .A1(n38308), .A2(n38743), .B1(n38306), .B2(n36303), .ZN(
        n8220) );
  OAI22_X1 U2465 ( .A1(n38309), .A2(n38750), .B1(n38306), .B2(n36304), .ZN(
        n8221) );
  OAI22_X1 U2466 ( .A1(n38309), .A2(n38757), .B1(n38306), .B2(n36305), .ZN(
        n8222) );
  OAI22_X1 U2467 ( .A1(n38309), .A2(n38764), .B1(n38306), .B2(n36306), .ZN(
        n8223) );
  OAI22_X1 U2468 ( .A1(n38309), .A2(n38771), .B1(n38306), .B2(n36307), .ZN(
        n8224) );
  OAI22_X1 U2469 ( .A1(n38309), .A2(n38778), .B1(n3831), .B2(n36308), .ZN(
        n8225) );
  OAI22_X1 U2470 ( .A1(n38310), .A2(n38785), .B1(n3831), .B2(n36309), .ZN(
        n8226) );
  OAI22_X1 U2471 ( .A1(n38310), .A2(n38792), .B1(n3831), .B2(n36310), .ZN(
        n8227) );
  OAI22_X1 U2472 ( .A1(n38310), .A2(n38799), .B1(n3831), .B2(n36311), .ZN(
        n8228) );
  OAI22_X1 U2473 ( .A1(n38310), .A2(n38806), .B1(n3831), .B2(n36312), .ZN(
        n8229) );
  OAI22_X1 U2474 ( .A1(n38310), .A2(n38813), .B1(n3831), .B2(n36313), .ZN(
        n8230) );
  OAI22_X1 U2475 ( .A1(n38311), .A2(n38820), .B1(n3831), .B2(n36314), .ZN(
        n8231) );
  OAI22_X1 U2476 ( .A1(n38311), .A2(n38827), .B1(n38306), .B2(n36315), .ZN(
        n8232) );
  OAI22_X1 U2477 ( .A1(n38311), .A2(n38834), .B1(n38306), .B2(n36316), .ZN(
        n8233) );
  OAI22_X1 U2478 ( .A1(n38311), .A2(n38841), .B1(n38306), .B2(n36317), .ZN(
        n8234) );
  OAI22_X1 U2479 ( .A1(n38319), .A2(n38680), .B1(n38318), .B2(n35566), .ZN(
        n8243) );
  OAI22_X1 U2480 ( .A1(n38319), .A2(n38687), .B1(n38318), .B2(n35568), .ZN(
        n8244) );
  OAI22_X1 U2481 ( .A1(n38319), .A2(n38694), .B1(n38318), .B2(n35570), .ZN(
        n8245) );
  OAI22_X1 U2482 ( .A1(n38319), .A2(n38701), .B1(n38318), .B2(n35572), .ZN(
        n8246) );
  OAI22_X1 U2483 ( .A1(n38319), .A2(n38708), .B1(n38318), .B2(n35574), .ZN(
        n8247) );
  OAI22_X1 U2484 ( .A1(n38320), .A2(n38715), .B1(n38318), .B2(n35576), .ZN(
        n8248) );
  OAI22_X1 U2485 ( .A1(n38320), .A2(n38722), .B1(n38318), .B2(n35578), .ZN(
        n8249) );
  OAI22_X1 U2486 ( .A1(n38320), .A2(n38729), .B1(n38318), .B2(n35580), .ZN(
        n8250) );
  OAI22_X1 U2487 ( .A1(n38320), .A2(n38736), .B1(n38318), .B2(n35582), .ZN(
        n8251) );
  OAI22_X1 U2488 ( .A1(n38320), .A2(n38743), .B1(n38318), .B2(n35584), .ZN(
        n8252) );
  OAI22_X1 U2489 ( .A1(n38321), .A2(n38750), .B1(n38318), .B2(n35586), .ZN(
        n8253) );
  OAI22_X1 U2490 ( .A1(n38321), .A2(n38757), .B1(n38318), .B2(n35588), .ZN(
        n8254) );
  OAI22_X1 U2491 ( .A1(n38321), .A2(n38764), .B1(n38318), .B2(n35590), .ZN(
        n8255) );
  OAI22_X1 U2492 ( .A1(n38321), .A2(n38771), .B1(n38318), .B2(n35592), .ZN(
        n8256) );
  OAI22_X1 U2493 ( .A1(n38321), .A2(n38778), .B1(n3796), .B2(n35594), .ZN(
        n8257) );
  OAI22_X1 U2494 ( .A1(n38322), .A2(n38785), .B1(n3796), .B2(n35596), .ZN(
        n8258) );
  OAI22_X1 U2495 ( .A1(n38322), .A2(n38792), .B1(n3796), .B2(n35598), .ZN(
        n8259) );
  OAI22_X1 U2496 ( .A1(n38322), .A2(n38799), .B1(n3796), .B2(n35600), .ZN(
        n8260) );
  OAI22_X1 U2497 ( .A1(n38322), .A2(n38806), .B1(n3796), .B2(n35602), .ZN(
        n8261) );
  OAI22_X1 U2498 ( .A1(n38322), .A2(n38813), .B1(n3796), .B2(n35604), .ZN(
        n8262) );
  OAI22_X1 U2499 ( .A1(n38323), .A2(n38820), .B1(n3796), .B2(n35606), .ZN(
        n8263) );
  OAI22_X1 U2500 ( .A1(n38323), .A2(n38827), .B1(n38318), .B2(n35608), .ZN(
        n8264) );
  OAI22_X1 U2501 ( .A1(n38323), .A2(n38834), .B1(n38318), .B2(n35610), .ZN(
        n8265) );
  OAI22_X1 U2502 ( .A1(n38323), .A2(n38841), .B1(n38318), .B2(n35612), .ZN(
        n8266) );
  OAI22_X1 U2503 ( .A1(n38340), .A2(n38679), .B1(n38339), .B2(n36638), .ZN(
        n8307) );
  OAI22_X1 U2504 ( .A1(n38340), .A2(n38686), .B1(n38339), .B2(n36640), .ZN(
        n8308) );
  OAI22_X1 U2505 ( .A1(n38340), .A2(n38693), .B1(n38339), .B2(n36642), .ZN(
        n8309) );
  OAI22_X1 U2506 ( .A1(n38340), .A2(n38700), .B1(n38339), .B2(n36644), .ZN(
        n8310) );
  OAI22_X1 U2507 ( .A1(n38340), .A2(n38707), .B1(n38339), .B2(n36646), .ZN(
        n8311) );
  OAI22_X1 U2508 ( .A1(n38341), .A2(n38714), .B1(n38339), .B2(n36648), .ZN(
        n8312) );
  OAI22_X1 U2509 ( .A1(n38341), .A2(n38721), .B1(n38339), .B2(n36650), .ZN(
        n8313) );
  OAI22_X1 U2510 ( .A1(n38341), .A2(n38728), .B1(n38339), .B2(n36652), .ZN(
        n8314) );
  OAI22_X1 U2511 ( .A1(n38341), .A2(n38735), .B1(n38339), .B2(n36654), .ZN(
        n8315) );
  OAI22_X1 U2512 ( .A1(n38341), .A2(n38742), .B1(n38339), .B2(n36656), .ZN(
        n8316) );
  OAI22_X1 U2513 ( .A1(n38342), .A2(n38749), .B1(n38339), .B2(n36658), .ZN(
        n8317) );
  OAI22_X1 U2514 ( .A1(n38342), .A2(n38756), .B1(n38339), .B2(n36660), .ZN(
        n8318) );
  OAI22_X1 U2515 ( .A1(n38342), .A2(n38763), .B1(n38339), .B2(n36662), .ZN(
        n8319) );
  OAI22_X1 U2516 ( .A1(n38342), .A2(n38770), .B1(n38339), .B2(n36664), .ZN(
        n8320) );
  OAI22_X1 U2517 ( .A1(n38342), .A2(n38777), .B1(n3726), .B2(n36666), .ZN(
        n8321) );
  OAI22_X1 U2518 ( .A1(n38343), .A2(n38784), .B1(n3726), .B2(n36668), .ZN(
        n8322) );
  OAI22_X1 U2519 ( .A1(n38343), .A2(n38791), .B1(n3726), .B2(n36670), .ZN(
        n8323) );
  OAI22_X1 U2520 ( .A1(n38343), .A2(n38798), .B1(n3726), .B2(n36672), .ZN(
        n8324) );
  OAI22_X1 U2521 ( .A1(n38343), .A2(n38805), .B1(n3726), .B2(n36674), .ZN(
        n8325) );
  OAI22_X1 U2522 ( .A1(n38343), .A2(n38812), .B1(n3726), .B2(n36676), .ZN(
        n8326) );
  OAI22_X1 U2523 ( .A1(n38344), .A2(n38819), .B1(n3726), .B2(n36678), .ZN(
        n8327) );
  OAI22_X1 U2524 ( .A1(n38344), .A2(n38826), .B1(n38339), .B2(n36680), .ZN(
        n8328) );
  OAI22_X1 U2525 ( .A1(n38344), .A2(n38833), .B1(n38339), .B2(n36682), .ZN(
        n8329) );
  OAI22_X1 U2526 ( .A1(n38344), .A2(n38840), .B1(n38339), .B2(n36684), .ZN(
        n8330) );
  OAI22_X1 U2527 ( .A1(n38361), .A2(n38679), .B1(n38360), .B2(n35928), .ZN(
        n8371) );
  OAI22_X1 U2528 ( .A1(n38361), .A2(n38686), .B1(n38360), .B2(n35932), .ZN(
        n8372) );
  OAI22_X1 U2529 ( .A1(n38361), .A2(n38693), .B1(n38360), .B2(n35936), .ZN(
        n8373) );
  OAI22_X1 U2530 ( .A1(n38361), .A2(n38700), .B1(n38360), .B2(n35940), .ZN(
        n8374) );
  OAI22_X1 U2531 ( .A1(n38361), .A2(n38707), .B1(n38360), .B2(n35944), .ZN(
        n8375) );
  OAI22_X1 U2532 ( .A1(n38362), .A2(n38714), .B1(n38360), .B2(n35948), .ZN(
        n8376) );
  OAI22_X1 U2533 ( .A1(n38362), .A2(n38721), .B1(n38360), .B2(n35952), .ZN(
        n8377) );
  OAI22_X1 U2534 ( .A1(n38362), .A2(n38728), .B1(n38360), .B2(n35956), .ZN(
        n8378) );
  OAI22_X1 U2535 ( .A1(n38362), .A2(n38735), .B1(n38360), .B2(n35960), .ZN(
        n8379) );
  OAI22_X1 U2536 ( .A1(n38362), .A2(n38742), .B1(n38360), .B2(n35964), .ZN(
        n8380) );
  OAI22_X1 U2537 ( .A1(n38363), .A2(n38749), .B1(n38360), .B2(n35968), .ZN(
        n8381) );
  OAI22_X1 U2538 ( .A1(n38363), .A2(n38756), .B1(n38360), .B2(n35972), .ZN(
        n8382) );
  OAI22_X1 U2539 ( .A1(n38363), .A2(n38763), .B1(n38360), .B2(n35976), .ZN(
        n8383) );
  OAI22_X1 U2540 ( .A1(n38363), .A2(n38770), .B1(n38360), .B2(n35980), .ZN(
        n8384) );
  OAI22_X1 U2541 ( .A1(n38363), .A2(n38777), .B1(n3656), .B2(n35984), .ZN(
        n8385) );
  OAI22_X1 U2542 ( .A1(n38364), .A2(n38784), .B1(n3656), .B2(n35988), .ZN(
        n8386) );
  OAI22_X1 U2543 ( .A1(n38364), .A2(n38791), .B1(n3656), .B2(n35992), .ZN(
        n8387) );
  OAI22_X1 U2544 ( .A1(n38364), .A2(n38798), .B1(n3656), .B2(n35996), .ZN(
        n8388) );
  OAI22_X1 U2545 ( .A1(n38364), .A2(n38805), .B1(n3656), .B2(n36000), .ZN(
        n8389) );
  OAI22_X1 U2546 ( .A1(n38364), .A2(n38812), .B1(n3656), .B2(n36004), .ZN(
        n8390) );
  OAI22_X1 U2547 ( .A1(n38365), .A2(n38819), .B1(n3656), .B2(n36008), .ZN(
        n8391) );
  OAI22_X1 U2548 ( .A1(n38365), .A2(n38826), .B1(n38360), .B2(n36012), .ZN(
        n8392) );
  OAI22_X1 U2549 ( .A1(n38365), .A2(n38833), .B1(n38360), .B2(n36016), .ZN(
        n8393) );
  OAI22_X1 U2550 ( .A1(n38365), .A2(n38840), .B1(n38360), .B2(n36020), .ZN(
        n8394) );
  OAI22_X1 U2551 ( .A1(n38373), .A2(n38679), .B1(n38372), .B2(n35518), .ZN(
        n8403) );
  OAI22_X1 U2552 ( .A1(n38373), .A2(n38686), .B1(n38372), .B2(n35520), .ZN(
        n8404) );
  OAI22_X1 U2553 ( .A1(n38373), .A2(n38693), .B1(n38372), .B2(n35522), .ZN(
        n8405) );
  OAI22_X1 U2554 ( .A1(n38373), .A2(n38700), .B1(n38372), .B2(n35524), .ZN(
        n8406) );
  OAI22_X1 U2555 ( .A1(n38373), .A2(n38707), .B1(n38372), .B2(n35526), .ZN(
        n8407) );
  OAI22_X1 U2556 ( .A1(n38374), .A2(n38714), .B1(n38372), .B2(n35528), .ZN(
        n8408) );
  OAI22_X1 U2557 ( .A1(n38374), .A2(n38721), .B1(n38372), .B2(n35530), .ZN(
        n8409) );
  OAI22_X1 U2558 ( .A1(n38374), .A2(n38728), .B1(n38372), .B2(n35532), .ZN(
        n8410) );
  OAI22_X1 U2559 ( .A1(n38374), .A2(n38735), .B1(n38372), .B2(n35534), .ZN(
        n8411) );
  OAI22_X1 U2560 ( .A1(n38374), .A2(n38742), .B1(n38372), .B2(n35536), .ZN(
        n8412) );
  OAI22_X1 U2561 ( .A1(n38375), .A2(n38749), .B1(n38372), .B2(n35538), .ZN(
        n8413) );
  OAI22_X1 U2562 ( .A1(n38375), .A2(n38756), .B1(n38372), .B2(n35540), .ZN(
        n8414) );
  OAI22_X1 U2563 ( .A1(n38375), .A2(n38763), .B1(n38372), .B2(n35542), .ZN(
        n8415) );
  OAI22_X1 U2564 ( .A1(n38375), .A2(n38770), .B1(n38372), .B2(n35544), .ZN(
        n8416) );
  OAI22_X1 U2565 ( .A1(n38375), .A2(n38777), .B1(n3621), .B2(n35546), .ZN(
        n8417) );
  OAI22_X1 U2566 ( .A1(n38376), .A2(n38784), .B1(n3621), .B2(n35548), .ZN(
        n8418) );
  OAI22_X1 U2567 ( .A1(n38376), .A2(n38791), .B1(n3621), .B2(n35550), .ZN(
        n8419) );
  OAI22_X1 U2568 ( .A1(n38376), .A2(n38798), .B1(n3621), .B2(n35552), .ZN(
        n8420) );
  OAI22_X1 U2569 ( .A1(n38376), .A2(n38805), .B1(n3621), .B2(n35554), .ZN(
        n8421) );
  OAI22_X1 U2570 ( .A1(n38376), .A2(n38812), .B1(n3621), .B2(n35556), .ZN(
        n8422) );
  OAI22_X1 U2571 ( .A1(n38377), .A2(n38819), .B1(n3621), .B2(n35558), .ZN(
        n8423) );
  OAI22_X1 U2572 ( .A1(n38377), .A2(n38826), .B1(n38372), .B2(n35560), .ZN(
        n8424) );
  OAI22_X1 U2573 ( .A1(n38377), .A2(n38833), .B1(n38372), .B2(n35562), .ZN(
        n8425) );
  OAI22_X1 U2574 ( .A1(n38377), .A2(n38840), .B1(n38372), .B2(n35564), .ZN(
        n8426) );
  OAI22_X1 U2575 ( .A1(n38394), .A2(n38679), .B1(n38393), .B2(n36591), .ZN(
        n8467) );
  OAI22_X1 U2576 ( .A1(n38394), .A2(n38686), .B1(n38393), .B2(n36593), .ZN(
        n8468) );
  OAI22_X1 U2577 ( .A1(n38394), .A2(n38693), .B1(n38393), .B2(n36595), .ZN(
        n8469) );
  OAI22_X1 U2578 ( .A1(n38394), .A2(n38700), .B1(n38393), .B2(n36597), .ZN(
        n8470) );
  OAI22_X1 U2579 ( .A1(n38394), .A2(n38707), .B1(n38393), .B2(n36599), .ZN(
        n8471) );
  OAI22_X1 U2580 ( .A1(n38395), .A2(n38714), .B1(n38393), .B2(n36601), .ZN(
        n8472) );
  OAI22_X1 U2581 ( .A1(n38395), .A2(n38721), .B1(n38393), .B2(n36603), .ZN(
        n8473) );
  OAI22_X1 U2582 ( .A1(n38395), .A2(n38728), .B1(n38393), .B2(n36605), .ZN(
        n8474) );
  OAI22_X1 U2583 ( .A1(n38395), .A2(n38735), .B1(n38393), .B2(n36607), .ZN(
        n8475) );
  OAI22_X1 U2584 ( .A1(n38395), .A2(n38742), .B1(n38393), .B2(n36609), .ZN(
        n8476) );
  OAI22_X1 U2585 ( .A1(n38396), .A2(n38749), .B1(n38393), .B2(n36611), .ZN(
        n8477) );
  OAI22_X1 U2586 ( .A1(n38396), .A2(n38756), .B1(n38393), .B2(n36613), .ZN(
        n8478) );
  OAI22_X1 U2587 ( .A1(n38396), .A2(n38763), .B1(n38393), .B2(n36615), .ZN(
        n8479) );
  OAI22_X1 U2588 ( .A1(n38396), .A2(n38770), .B1(n38393), .B2(n36617), .ZN(
        n8480) );
  OAI22_X1 U2589 ( .A1(n38396), .A2(n38777), .B1(n3551), .B2(n36619), .ZN(
        n8481) );
  OAI22_X1 U2590 ( .A1(n38397), .A2(n38784), .B1(n3551), .B2(n36621), .ZN(
        n8482) );
  OAI22_X1 U2591 ( .A1(n38397), .A2(n38791), .B1(n3551), .B2(n36623), .ZN(
        n8483) );
  OAI22_X1 U2592 ( .A1(n38397), .A2(n38798), .B1(n3551), .B2(n36625), .ZN(
        n8484) );
  OAI22_X1 U2593 ( .A1(n38397), .A2(n38805), .B1(n3551), .B2(n36627), .ZN(
        n8485) );
  OAI22_X1 U2594 ( .A1(n38397), .A2(n38812), .B1(n3551), .B2(n36629), .ZN(
        n8486) );
  OAI22_X1 U2595 ( .A1(n38398), .A2(n38819), .B1(n3551), .B2(n36631), .ZN(
        n8487) );
  OAI22_X1 U2596 ( .A1(n38398), .A2(n38826), .B1(n38393), .B2(n36633), .ZN(
        n8488) );
  OAI22_X1 U2597 ( .A1(n38398), .A2(n38833), .B1(n38393), .B2(n36635), .ZN(
        n8489) );
  OAI22_X1 U2598 ( .A1(n38398), .A2(n38840), .B1(n38393), .B2(n36637), .ZN(
        n8490) );
  OAI22_X1 U2599 ( .A1(n38415), .A2(n38679), .B1(n38414), .B2(n36127), .ZN(
        n8531) );
  OAI22_X1 U2600 ( .A1(n38415), .A2(n38686), .B1(n38414), .B2(n36129), .ZN(
        n8532) );
  OAI22_X1 U2601 ( .A1(n38415), .A2(n38693), .B1(n38414), .B2(n36131), .ZN(
        n8533) );
  OAI22_X1 U2602 ( .A1(n38415), .A2(n38700), .B1(n38414), .B2(n36133), .ZN(
        n8534) );
  OAI22_X1 U2603 ( .A1(n38415), .A2(n38707), .B1(n38414), .B2(n36135), .ZN(
        n8535) );
  OAI22_X1 U2604 ( .A1(n38416), .A2(n38714), .B1(n38414), .B2(n36137), .ZN(
        n8536) );
  OAI22_X1 U2605 ( .A1(n38416), .A2(n38721), .B1(n38414), .B2(n36139), .ZN(
        n8537) );
  OAI22_X1 U2606 ( .A1(n38416), .A2(n38728), .B1(n38414), .B2(n36141), .ZN(
        n8538) );
  OAI22_X1 U2607 ( .A1(n38416), .A2(n38735), .B1(n38414), .B2(n36143), .ZN(
        n8539) );
  OAI22_X1 U2608 ( .A1(n38416), .A2(n38742), .B1(n38414), .B2(n36145), .ZN(
        n8540) );
  OAI22_X1 U2609 ( .A1(n38417), .A2(n38749), .B1(n38414), .B2(n36147), .ZN(
        n8541) );
  OAI22_X1 U2610 ( .A1(n38417), .A2(n38756), .B1(n38414), .B2(n36149), .ZN(
        n8542) );
  OAI22_X1 U2611 ( .A1(n38417), .A2(n38763), .B1(n38414), .B2(n36151), .ZN(
        n8543) );
  OAI22_X1 U2612 ( .A1(n38417), .A2(n38770), .B1(n38414), .B2(n36153), .ZN(
        n8544) );
  OAI22_X1 U2613 ( .A1(n38417), .A2(n38777), .B1(n3481), .B2(n36155), .ZN(
        n8545) );
  OAI22_X1 U2614 ( .A1(n38418), .A2(n38784), .B1(n3481), .B2(n36157), .ZN(
        n8546) );
  OAI22_X1 U2615 ( .A1(n38418), .A2(n38791), .B1(n3481), .B2(n36159), .ZN(
        n8547) );
  OAI22_X1 U2616 ( .A1(n38418), .A2(n38798), .B1(n3481), .B2(n36161), .ZN(
        n8548) );
  OAI22_X1 U2617 ( .A1(n38418), .A2(n38805), .B1(n3481), .B2(n36163), .ZN(
        n8549) );
  OAI22_X1 U2618 ( .A1(n38418), .A2(n38812), .B1(n3481), .B2(n36165), .ZN(
        n8550) );
  OAI22_X1 U2619 ( .A1(n38419), .A2(n38819), .B1(n3481), .B2(n36167), .ZN(
        n8551) );
  OAI22_X1 U2620 ( .A1(n38419), .A2(n38826), .B1(n38414), .B2(n36169), .ZN(
        n8552) );
  OAI22_X1 U2621 ( .A1(n38419), .A2(n38833), .B1(n38414), .B2(n36171), .ZN(
        n8553) );
  OAI22_X1 U2622 ( .A1(n38419), .A2(n38840), .B1(n38414), .B2(n36173), .ZN(
        n8554) );
  OAI22_X1 U2623 ( .A1(n38427), .A2(n38679), .B1(n38426), .B2(n35417), .ZN(
        n8563) );
  OAI22_X1 U2624 ( .A1(n38427), .A2(n38686), .B1(n38426), .B2(n35421), .ZN(
        n8564) );
  OAI22_X1 U2625 ( .A1(n38427), .A2(n38693), .B1(n38426), .B2(n35425), .ZN(
        n8565) );
  OAI22_X1 U2626 ( .A1(n38427), .A2(n38700), .B1(n38426), .B2(n35429), .ZN(
        n8566) );
  OAI22_X1 U2627 ( .A1(n38427), .A2(n38707), .B1(n38426), .B2(n35433), .ZN(
        n8567) );
  OAI22_X1 U2628 ( .A1(n38428), .A2(n38714), .B1(n38426), .B2(n35437), .ZN(
        n8568) );
  OAI22_X1 U2629 ( .A1(n38428), .A2(n38721), .B1(n38426), .B2(n35441), .ZN(
        n8569) );
  OAI22_X1 U2630 ( .A1(n38428), .A2(n38728), .B1(n38426), .B2(n35445), .ZN(
        n8570) );
  OAI22_X1 U2631 ( .A1(n38428), .A2(n38735), .B1(n38426), .B2(n35449), .ZN(
        n8571) );
  OAI22_X1 U2632 ( .A1(n38428), .A2(n38742), .B1(n38426), .B2(n35453), .ZN(
        n8572) );
  OAI22_X1 U2633 ( .A1(n38429), .A2(n38749), .B1(n38426), .B2(n35457), .ZN(
        n8573) );
  OAI22_X1 U2634 ( .A1(n38429), .A2(n38756), .B1(n38426), .B2(n35461), .ZN(
        n8574) );
  OAI22_X1 U2635 ( .A1(n38429), .A2(n38763), .B1(n38426), .B2(n35465), .ZN(
        n8575) );
  OAI22_X1 U2636 ( .A1(n38429), .A2(n38770), .B1(n38426), .B2(n35469), .ZN(
        n8576) );
  OAI22_X1 U2637 ( .A1(n38429), .A2(n38777), .B1(n3446), .B2(n35473), .ZN(
        n8577) );
  OAI22_X1 U2638 ( .A1(n38430), .A2(n38784), .B1(n3446), .B2(n35477), .ZN(
        n8578) );
  OAI22_X1 U2639 ( .A1(n38430), .A2(n38791), .B1(n3446), .B2(n35481), .ZN(
        n8579) );
  OAI22_X1 U2640 ( .A1(n38430), .A2(n38798), .B1(n3446), .B2(n35485), .ZN(
        n8580) );
  OAI22_X1 U2641 ( .A1(n38430), .A2(n38805), .B1(n3446), .B2(n35489), .ZN(
        n8581) );
  OAI22_X1 U2642 ( .A1(n38430), .A2(n38812), .B1(n3446), .B2(n35493), .ZN(
        n8582) );
  OAI22_X1 U2643 ( .A1(n38431), .A2(n38819), .B1(n3446), .B2(n35497), .ZN(
        n8583) );
  OAI22_X1 U2644 ( .A1(n38431), .A2(n38826), .B1(n38426), .B2(n35501), .ZN(
        n8584) );
  OAI22_X1 U2645 ( .A1(n38431), .A2(n38833), .B1(n38426), .B2(n35505), .ZN(
        n8585) );
  OAI22_X1 U2646 ( .A1(n38431), .A2(n38840), .B1(n38426), .B2(n35509), .ZN(
        n8586) );
  OAI22_X1 U2647 ( .A1(n38448), .A2(n38679), .B1(n38447), .B2(n36543), .ZN(
        n8627) );
  OAI22_X1 U2648 ( .A1(n38448), .A2(n38686), .B1(n38447), .B2(n36545), .ZN(
        n8628) );
  OAI22_X1 U2649 ( .A1(n38448), .A2(n38693), .B1(n38447), .B2(n36547), .ZN(
        n8629) );
  OAI22_X1 U2650 ( .A1(n38448), .A2(n38700), .B1(n38447), .B2(n36549), .ZN(
        n8630) );
  OAI22_X1 U2651 ( .A1(n38448), .A2(n38707), .B1(n38447), .B2(n36551), .ZN(
        n8631) );
  OAI22_X1 U2652 ( .A1(n38449), .A2(n38714), .B1(n38447), .B2(n36553), .ZN(
        n8632) );
  OAI22_X1 U2653 ( .A1(n38449), .A2(n38721), .B1(n38447), .B2(n36555), .ZN(
        n8633) );
  OAI22_X1 U2654 ( .A1(n38449), .A2(n38728), .B1(n38447), .B2(n36557), .ZN(
        n8634) );
  OAI22_X1 U2655 ( .A1(n38449), .A2(n38735), .B1(n38447), .B2(n36559), .ZN(
        n8635) );
  OAI22_X1 U2656 ( .A1(n38449), .A2(n38742), .B1(n38447), .B2(n36561), .ZN(
        n8636) );
  OAI22_X1 U2657 ( .A1(n38450), .A2(n38749), .B1(n38447), .B2(n36563), .ZN(
        n8637) );
  OAI22_X1 U2658 ( .A1(n38450), .A2(n38756), .B1(n38447), .B2(n36565), .ZN(
        n8638) );
  OAI22_X1 U2659 ( .A1(n38450), .A2(n38763), .B1(n38447), .B2(n36567), .ZN(
        n8639) );
  OAI22_X1 U2660 ( .A1(n38450), .A2(n38770), .B1(n38447), .B2(n36569), .ZN(
        n8640) );
  OAI22_X1 U2661 ( .A1(n38450), .A2(n38777), .B1(n3376), .B2(n36571), .ZN(
        n8641) );
  OAI22_X1 U2662 ( .A1(n38451), .A2(n38784), .B1(n3376), .B2(n36573), .ZN(
        n8642) );
  OAI22_X1 U2663 ( .A1(n38451), .A2(n38791), .B1(n3376), .B2(n36575), .ZN(
        n8643) );
  OAI22_X1 U2664 ( .A1(n38451), .A2(n38798), .B1(n3376), .B2(n36577), .ZN(
        n8644) );
  OAI22_X1 U2665 ( .A1(n38451), .A2(n38805), .B1(n3376), .B2(n36579), .ZN(
        n8645) );
  OAI22_X1 U2666 ( .A1(n38451), .A2(n38812), .B1(n3376), .B2(n36581), .ZN(
        n8646) );
  OAI22_X1 U2667 ( .A1(n38452), .A2(n38819), .B1(n3376), .B2(n36583), .ZN(
        n8647) );
  OAI22_X1 U2668 ( .A1(n38452), .A2(n38826), .B1(n38447), .B2(n36585), .ZN(
        n8648) );
  OAI22_X1 U2669 ( .A1(n38452), .A2(n38833), .B1(n38447), .B2(n36587), .ZN(
        n8649) );
  OAI22_X1 U2670 ( .A1(n38452), .A2(n38840), .B1(n38447), .B2(n36589), .ZN(
        n8650) );
  OAI22_X1 U2671 ( .A1(n38469), .A2(n38678), .B1(n38468), .B2(n35782), .ZN(
        n8691) );
  OAI22_X1 U2672 ( .A1(n38469), .A2(n38685), .B1(n38468), .B2(n35783), .ZN(
        n8692) );
  OAI22_X1 U2673 ( .A1(n38469), .A2(n38692), .B1(n38468), .B2(n35784), .ZN(
        n8693) );
  OAI22_X1 U2674 ( .A1(n38469), .A2(n38699), .B1(n38468), .B2(n35785), .ZN(
        n8694) );
  OAI22_X1 U2675 ( .A1(n38469), .A2(n38706), .B1(n38468), .B2(n35786), .ZN(
        n8695) );
  OAI22_X1 U2676 ( .A1(n38470), .A2(n38713), .B1(n38468), .B2(n35787), .ZN(
        n8696) );
  OAI22_X1 U2677 ( .A1(n38470), .A2(n38720), .B1(n38468), .B2(n35788), .ZN(
        n8697) );
  OAI22_X1 U2678 ( .A1(n38470), .A2(n38727), .B1(n38468), .B2(n35789), .ZN(
        n8698) );
  OAI22_X1 U2679 ( .A1(n38470), .A2(n38734), .B1(n38468), .B2(n35790), .ZN(
        n8699) );
  OAI22_X1 U2680 ( .A1(n38470), .A2(n38741), .B1(n38468), .B2(n35791), .ZN(
        n8700) );
  OAI22_X1 U2681 ( .A1(n38471), .A2(n38748), .B1(n38468), .B2(n35792), .ZN(
        n8701) );
  OAI22_X1 U2682 ( .A1(n38471), .A2(n38755), .B1(n38468), .B2(n35793), .ZN(
        n8702) );
  OAI22_X1 U2683 ( .A1(n38471), .A2(n38762), .B1(n38468), .B2(n35794), .ZN(
        n8703) );
  OAI22_X1 U2684 ( .A1(n38471), .A2(n38769), .B1(n38468), .B2(n35795), .ZN(
        n8704) );
  OAI22_X1 U2685 ( .A1(n38471), .A2(n38776), .B1(n3306), .B2(n35796), .ZN(
        n8705) );
  OAI22_X1 U2686 ( .A1(n38472), .A2(n38783), .B1(n3306), .B2(n35797), .ZN(
        n8706) );
  OAI22_X1 U2687 ( .A1(n38472), .A2(n38790), .B1(n3306), .B2(n35798), .ZN(
        n8707) );
  OAI22_X1 U2688 ( .A1(n38472), .A2(n38797), .B1(n3306), .B2(n35799), .ZN(
        n8708) );
  OAI22_X1 U2689 ( .A1(n38472), .A2(n38804), .B1(n3306), .B2(n35800), .ZN(
        n8709) );
  OAI22_X1 U2690 ( .A1(n38472), .A2(n38811), .B1(n3306), .B2(n35801), .ZN(
        n8710) );
  OAI22_X1 U2691 ( .A1(n38473), .A2(n38818), .B1(n3306), .B2(n35802), .ZN(
        n8711) );
  OAI22_X1 U2692 ( .A1(n38473), .A2(n38825), .B1(n38468), .B2(n35803), .ZN(
        n8712) );
  OAI22_X1 U2693 ( .A1(n38473), .A2(n38832), .B1(n38468), .B2(n35804), .ZN(
        n8713) );
  OAI22_X1 U2694 ( .A1(n38473), .A2(n38839), .B1(n38468), .B2(n35805), .ZN(
        n8714) );
  OAI22_X1 U2695 ( .A1(n38487), .A2(n38678), .B1(n38486), .B2(n35270), .ZN(
        n8723) );
  OAI22_X1 U2696 ( .A1(n38487), .A2(n38685), .B1(n38486), .B2(n35271), .ZN(
        n8724) );
  OAI22_X1 U2697 ( .A1(n38487), .A2(n38692), .B1(n38486), .B2(n35272), .ZN(
        n8725) );
  OAI22_X1 U2698 ( .A1(n38487), .A2(n38699), .B1(n38486), .B2(n35273), .ZN(
        n8726) );
  OAI22_X1 U2699 ( .A1(n38487), .A2(n38706), .B1(n38486), .B2(n35274), .ZN(
        n8727) );
  OAI22_X1 U2700 ( .A1(n38488), .A2(n38713), .B1(n38486), .B2(n35275), .ZN(
        n8728) );
  OAI22_X1 U2701 ( .A1(n38488), .A2(n38720), .B1(n38486), .B2(n35276), .ZN(
        n8729) );
  OAI22_X1 U2702 ( .A1(n38488), .A2(n38727), .B1(n38486), .B2(n35277), .ZN(
        n8730) );
  OAI22_X1 U2703 ( .A1(n38488), .A2(n38734), .B1(n38486), .B2(n35278), .ZN(
        n8731) );
  OAI22_X1 U2704 ( .A1(n38488), .A2(n38741), .B1(n38486), .B2(n35279), .ZN(
        n8732) );
  OAI22_X1 U2705 ( .A1(n38489), .A2(n38748), .B1(n38486), .B2(n35280), .ZN(
        n8733) );
  OAI22_X1 U2706 ( .A1(n38489), .A2(n38755), .B1(n38486), .B2(n35281), .ZN(
        n8734) );
  OAI22_X1 U2707 ( .A1(n38489), .A2(n38762), .B1(n38486), .B2(n35282), .ZN(
        n8735) );
  OAI22_X1 U2708 ( .A1(n38489), .A2(n38769), .B1(n38486), .B2(n35283), .ZN(
        n8736) );
  OAI22_X1 U2709 ( .A1(n38489), .A2(n38776), .B1(n3270), .B2(n35284), .ZN(
        n8737) );
  OAI22_X1 U2710 ( .A1(n38490), .A2(n38783), .B1(n3270), .B2(n35285), .ZN(
        n8738) );
  OAI22_X1 U2711 ( .A1(n38490), .A2(n38790), .B1(n3270), .B2(n35286), .ZN(
        n8739) );
  OAI22_X1 U2712 ( .A1(n38490), .A2(n38797), .B1(n3270), .B2(n35287), .ZN(
        n8740) );
  OAI22_X1 U2713 ( .A1(n38490), .A2(n38804), .B1(n3270), .B2(n35288), .ZN(
        n8741) );
  OAI22_X1 U2714 ( .A1(n38490), .A2(n38811), .B1(n3270), .B2(n35289), .ZN(
        n8742) );
  OAI22_X1 U2715 ( .A1(n38491), .A2(n38818), .B1(n3270), .B2(n35290), .ZN(
        n8743) );
  OAI22_X1 U2716 ( .A1(n38491), .A2(n38825), .B1(n38486), .B2(n35291), .ZN(
        n8744) );
  OAI22_X1 U2717 ( .A1(n38491), .A2(n38832), .B1(n38486), .B2(n35292), .ZN(
        n8745) );
  OAI22_X1 U2718 ( .A1(n38491), .A2(n38839), .B1(n38486), .B2(n35293), .ZN(
        n8746) );
  OAI22_X1 U2719 ( .A1(n38511), .A2(n38678), .B1(n38510), .B2(n35294), .ZN(
        n8787) );
  OAI22_X1 U2720 ( .A1(n38511), .A2(n38685), .B1(n38510), .B2(n35295), .ZN(
        n8788) );
  OAI22_X1 U2721 ( .A1(n38511), .A2(n38692), .B1(n38510), .B2(n35296), .ZN(
        n8789) );
  OAI22_X1 U2722 ( .A1(n38511), .A2(n38699), .B1(n38510), .B2(n35297), .ZN(
        n8790) );
  OAI22_X1 U2723 ( .A1(n38511), .A2(n38706), .B1(n38510), .B2(n35298), .ZN(
        n8791) );
  OAI22_X1 U2724 ( .A1(n38512), .A2(n38713), .B1(n38510), .B2(n35299), .ZN(
        n8792) );
  OAI22_X1 U2725 ( .A1(n38512), .A2(n38720), .B1(n38510), .B2(n35300), .ZN(
        n8793) );
  OAI22_X1 U2726 ( .A1(n38512), .A2(n38727), .B1(n38510), .B2(n35301), .ZN(
        n8794) );
  OAI22_X1 U2727 ( .A1(n38512), .A2(n38734), .B1(n38510), .B2(n35302), .ZN(
        n8795) );
  OAI22_X1 U2728 ( .A1(n38512), .A2(n38741), .B1(n38510), .B2(n35303), .ZN(
        n8796) );
  OAI22_X1 U2729 ( .A1(n38513), .A2(n38748), .B1(n38510), .B2(n35304), .ZN(
        n8797) );
  OAI22_X1 U2730 ( .A1(n38513), .A2(n38755), .B1(n38510), .B2(n35305), .ZN(
        n8798) );
  OAI22_X1 U2731 ( .A1(n38513), .A2(n38762), .B1(n3200), .B2(n35306), .ZN(
        n8799) );
  OAI22_X1 U2732 ( .A1(n38513), .A2(n38769), .B1(n3200), .B2(n35307), .ZN(
        n8800) );
  OAI22_X1 U2733 ( .A1(n38513), .A2(n38776), .B1(n3200), .B2(n35308), .ZN(
        n8801) );
  OAI22_X1 U2734 ( .A1(n38514), .A2(n38783), .B1(n3200), .B2(n35309), .ZN(
        n8802) );
  OAI22_X1 U2735 ( .A1(n38514), .A2(n38790), .B1(n3200), .B2(n35310), .ZN(
        n8803) );
  OAI22_X1 U2736 ( .A1(n38514), .A2(n38797), .B1(n3200), .B2(n35311), .ZN(
        n8804) );
  OAI22_X1 U2737 ( .A1(n38514), .A2(n38804), .B1(n3200), .B2(n35312), .ZN(
        n8805) );
  OAI22_X1 U2738 ( .A1(n38514), .A2(n38811), .B1(n3200), .B2(n35313), .ZN(
        n8806) );
  OAI22_X1 U2739 ( .A1(n38515), .A2(n38818), .B1(n3200), .B2(n35314), .ZN(
        n8807) );
  OAI22_X1 U2740 ( .A1(n38515), .A2(n38825), .B1(n38510), .B2(n35315), .ZN(
        n8808) );
  OAI22_X1 U2741 ( .A1(n38515), .A2(n38832), .B1(n38510), .B2(n35316), .ZN(
        n8809) );
  OAI22_X1 U2742 ( .A1(n38515), .A2(n38839), .B1(n38510), .B2(n35317), .ZN(
        n8810) );
  OAI22_X1 U2743 ( .A1(n38523), .A2(n38678), .B1(n38522), .B2(n36318), .ZN(
        n8819) );
  OAI22_X1 U2744 ( .A1(n38523), .A2(n38685), .B1(n38522), .B2(n36319), .ZN(
        n8820) );
  OAI22_X1 U2745 ( .A1(n38523), .A2(n38692), .B1(n38522), .B2(n36320), .ZN(
        n8821) );
  OAI22_X1 U2746 ( .A1(n38523), .A2(n38699), .B1(n38522), .B2(n36321), .ZN(
        n8822) );
  OAI22_X1 U2747 ( .A1(n38523), .A2(n38706), .B1(n38522), .B2(n36322), .ZN(
        n8823) );
  OAI22_X1 U2748 ( .A1(n38524), .A2(n38713), .B1(n38522), .B2(n36323), .ZN(
        n8824) );
  OAI22_X1 U2749 ( .A1(n38524), .A2(n38720), .B1(n38522), .B2(n36324), .ZN(
        n8825) );
  OAI22_X1 U2750 ( .A1(n38524), .A2(n38727), .B1(n38522), .B2(n36325), .ZN(
        n8826) );
  OAI22_X1 U2751 ( .A1(n38524), .A2(n38734), .B1(n38522), .B2(n36326), .ZN(
        n8827) );
  OAI22_X1 U2752 ( .A1(n38524), .A2(n38741), .B1(n38522), .B2(n36327), .ZN(
        n8828) );
  OAI22_X1 U2753 ( .A1(n38525), .A2(n38748), .B1(n38522), .B2(n36328), .ZN(
        n8829) );
  OAI22_X1 U2754 ( .A1(n38525), .A2(n38755), .B1(n38522), .B2(n36329), .ZN(
        n8830) );
  OAI22_X1 U2755 ( .A1(n38525), .A2(n38762), .B1(n3165), .B2(n36330), .ZN(
        n8831) );
  OAI22_X1 U2756 ( .A1(n38525), .A2(n38769), .B1(n3165), .B2(n36331), .ZN(
        n8832) );
  OAI22_X1 U2757 ( .A1(n38525), .A2(n38776), .B1(n3165), .B2(n36332), .ZN(
        n8833) );
  OAI22_X1 U2758 ( .A1(n38526), .A2(n38783), .B1(n3165), .B2(n36333), .ZN(
        n8834) );
  OAI22_X1 U2759 ( .A1(n38526), .A2(n38790), .B1(n3165), .B2(n36334), .ZN(
        n8835) );
  OAI22_X1 U2760 ( .A1(n38526), .A2(n38797), .B1(n3165), .B2(n36335), .ZN(
        n8836) );
  OAI22_X1 U2761 ( .A1(n38526), .A2(n38804), .B1(n3165), .B2(n36336), .ZN(
        n8837) );
  OAI22_X1 U2762 ( .A1(n38526), .A2(n38811), .B1(n3165), .B2(n36337), .ZN(
        n8838) );
  OAI22_X1 U2763 ( .A1(n38527), .A2(n38818), .B1(n3165), .B2(n36338), .ZN(
        n8839) );
  OAI22_X1 U2764 ( .A1(n38527), .A2(n38825), .B1(n38522), .B2(n36339), .ZN(
        n8840) );
  OAI22_X1 U2765 ( .A1(n38527), .A2(n38832), .B1(n38522), .B2(n36340), .ZN(
        n8841) );
  OAI22_X1 U2766 ( .A1(n38527), .A2(n38839), .B1(n38522), .B2(n36341), .ZN(
        n8842) );
  OAI22_X1 U2767 ( .A1(n38535), .A2(n38678), .B1(n38534), .B2(n35806), .ZN(
        n8851) );
  OAI22_X1 U2768 ( .A1(n38535), .A2(n38685), .B1(n38534), .B2(n35807), .ZN(
        n8852) );
  OAI22_X1 U2769 ( .A1(n38535), .A2(n38692), .B1(n38534), .B2(n35808), .ZN(
        n8853) );
  OAI22_X1 U2770 ( .A1(n38535), .A2(n38699), .B1(n38534), .B2(n35809), .ZN(
        n8854) );
  OAI22_X1 U2771 ( .A1(n38535), .A2(n38706), .B1(n38534), .B2(n35810), .ZN(
        n8855) );
  OAI22_X1 U2772 ( .A1(n38536), .A2(n38713), .B1(n38534), .B2(n35811), .ZN(
        n8856) );
  OAI22_X1 U2773 ( .A1(n38536), .A2(n38720), .B1(n38534), .B2(n35812), .ZN(
        n8857) );
  OAI22_X1 U2774 ( .A1(n38536), .A2(n38727), .B1(n38534), .B2(n35813), .ZN(
        n8858) );
  OAI22_X1 U2775 ( .A1(n38536), .A2(n38734), .B1(n38534), .B2(n35814), .ZN(
        n8859) );
  OAI22_X1 U2776 ( .A1(n38536), .A2(n38741), .B1(n38534), .B2(n35815), .ZN(
        n8860) );
  OAI22_X1 U2777 ( .A1(n38537), .A2(n38748), .B1(n38534), .B2(n35816), .ZN(
        n8861) );
  OAI22_X1 U2778 ( .A1(n38537), .A2(n38755), .B1(n38534), .B2(n35817), .ZN(
        n8862) );
  OAI22_X1 U2779 ( .A1(n38537), .A2(n38762), .B1(n3130), .B2(n35818), .ZN(
        n8863) );
  OAI22_X1 U2780 ( .A1(n38537), .A2(n38769), .B1(n3130), .B2(n35819), .ZN(
        n8864) );
  OAI22_X1 U2781 ( .A1(n38537), .A2(n38776), .B1(n3130), .B2(n35820), .ZN(
        n8865) );
  OAI22_X1 U2782 ( .A1(n38538), .A2(n38783), .B1(n3130), .B2(n35821), .ZN(
        n8866) );
  OAI22_X1 U2783 ( .A1(n38538), .A2(n38790), .B1(n3130), .B2(n35822), .ZN(
        n8867) );
  OAI22_X1 U2784 ( .A1(n38538), .A2(n38797), .B1(n3130), .B2(n35823), .ZN(
        n8868) );
  OAI22_X1 U2785 ( .A1(n38538), .A2(n38804), .B1(n3130), .B2(n35824), .ZN(
        n8869) );
  OAI22_X1 U2786 ( .A1(n38538), .A2(n38811), .B1(n3130), .B2(n35825), .ZN(
        n8870) );
  OAI22_X1 U2787 ( .A1(n38539), .A2(n38818), .B1(n3130), .B2(n35826), .ZN(
        n8871) );
  OAI22_X1 U2788 ( .A1(n38539), .A2(n38825), .B1(n38534), .B2(n35827), .ZN(
        n8872) );
  OAI22_X1 U2789 ( .A1(n38539), .A2(n38832), .B1(n38534), .B2(n35828), .ZN(
        n8873) );
  OAI22_X1 U2790 ( .A1(n38539), .A2(n38839), .B1(n38534), .B2(n35829), .ZN(
        n8874) );
  OAI22_X1 U2791 ( .A1(n38571), .A2(n38678), .B1(n38570), .B2(n35415), .ZN(
        n8947) );
  OAI22_X1 U2792 ( .A1(n38571), .A2(n38685), .B1(n38570), .B2(n35419), .ZN(
        n8948) );
  OAI22_X1 U2793 ( .A1(n38571), .A2(n38692), .B1(n38570), .B2(n35423), .ZN(
        n8949) );
  OAI22_X1 U2794 ( .A1(n38571), .A2(n38699), .B1(n38570), .B2(n35427), .ZN(
        n8950) );
  OAI22_X1 U2795 ( .A1(n38571), .A2(n38706), .B1(n38570), .B2(n35431), .ZN(
        n8951) );
  OAI22_X1 U2796 ( .A1(n38572), .A2(n38713), .B1(n38570), .B2(n35435), .ZN(
        n8952) );
  OAI22_X1 U2797 ( .A1(n38572), .A2(n38720), .B1(n38570), .B2(n35439), .ZN(
        n8953) );
  OAI22_X1 U2798 ( .A1(n38572), .A2(n38727), .B1(n38570), .B2(n35443), .ZN(
        n8954) );
  OAI22_X1 U2799 ( .A1(n38572), .A2(n38734), .B1(n38570), .B2(n35447), .ZN(
        n8955) );
  OAI22_X1 U2800 ( .A1(n38572), .A2(n38741), .B1(n38570), .B2(n35451), .ZN(
        n8956) );
  OAI22_X1 U2801 ( .A1(n38573), .A2(n38748), .B1(n38570), .B2(n35455), .ZN(
        n8957) );
  OAI22_X1 U2802 ( .A1(n38573), .A2(n38755), .B1(n38570), .B2(n35459), .ZN(
        n8958) );
  OAI22_X1 U2803 ( .A1(n38573), .A2(n38762), .B1(n3025), .B2(n35463), .ZN(
        n8959) );
  OAI22_X1 U2804 ( .A1(n38573), .A2(n38769), .B1(n3025), .B2(n35467), .ZN(
        n8960) );
  OAI22_X1 U2805 ( .A1(n38573), .A2(n38776), .B1(n3025), .B2(n35471), .ZN(
        n8961) );
  OAI22_X1 U2806 ( .A1(n38574), .A2(n38783), .B1(n3025), .B2(n35475), .ZN(
        n8962) );
  OAI22_X1 U2807 ( .A1(n38574), .A2(n38790), .B1(n3025), .B2(n35479), .ZN(
        n8963) );
  OAI22_X1 U2808 ( .A1(n38574), .A2(n38797), .B1(n3025), .B2(n35483), .ZN(
        n8964) );
  OAI22_X1 U2809 ( .A1(n38574), .A2(n38804), .B1(n3025), .B2(n35487), .ZN(
        n8965) );
  OAI22_X1 U2810 ( .A1(n38574), .A2(n38811), .B1(n3025), .B2(n35491), .ZN(
        n8966) );
  OAI22_X1 U2811 ( .A1(n38575), .A2(n38818), .B1(n3025), .B2(n35495), .ZN(
        n8967) );
  OAI22_X1 U2812 ( .A1(n38575), .A2(n38825), .B1(n38570), .B2(n35499), .ZN(
        n8968) );
  OAI22_X1 U2813 ( .A1(n38575), .A2(n38832), .B1(n38570), .B2(n35503), .ZN(
        n8969) );
  OAI22_X1 U2814 ( .A1(n38575), .A2(n38839), .B1(n38570), .B2(n35507), .ZN(
        n8970) );
  OAI22_X1 U2815 ( .A1(n38583), .A2(n38678), .B1(n38582), .B2(n36439), .ZN(
        n8979) );
  OAI22_X1 U2816 ( .A1(n38583), .A2(n38685), .B1(n38582), .B2(n36443), .ZN(
        n8980) );
  OAI22_X1 U2817 ( .A1(n38583), .A2(n38692), .B1(n38582), .B2(n36447), .ZN(
        n8981) );
  OAI22_X1 U2818 ( .A1(n38583), .A2(n38699), .B1(n38582), .B2(n36451), .ZN(
        n8982) );
  OAI22_X1 U2819 ( .A1(n38583), .A2(n38706), .B1(n38582), .B2(n36455), .ZN(
        n8983) );
  OAI22_X1 U2820 ( .A1(n38584), .A2(n38713), .B1(n38582), .B2(n36459), .ZN(
        n8984) );
  OAI22_X1 U2821 ( .A1(n38584), .A2(n38720), .B1(n38582), .B2(n36463), .ZN(
        n8985) );
  OAI22_X1 U2822 ( .A1(n38584), .A2(n38727), .B1(n38582), .B2(n36467), .ZN(
        n8986) );
  OAI22_X1 U2823 ( .A1(n38584), .A2(n38734), .B1(n38582), .B2(n36471), .ZN(
        n8987) );
  OAI22_X1 U2824 ( .A1(n38584), .A2(n38741), .B1(n38582), .B2(n36475), .ZN(
        n8988) );
  OAI22_X1 U2825 ( .A1(n38585), .A2(n38748), .B1(n38582), .B2(n36479), .ZN(
        n8989) );
  OAI22_X1 U2826 ( .A1(n38585), .A2(n38755), .B1(n38582), .B2(n36483), .ZN(
        n8990) );
  OAI22_X1 U2827 ( .A1(n38585), .A2(n38762), .B1(n2990), .B2(n36487), .ZN(
        n8991) );
  OAI22_X1 U2828 ( .A1(n38585), .A2(n38769), .B1(n2990), .B2(n36491), .ZN(
        n8992) );
  OAI22_X1 U2829 ( .A1(n38585), .A2(n38776), .B1(n2990), .B2(n36495), .ZN(
        n8993) );
  OAI22_X1 U2830 ( .A1(n38586), .A2(n38783), .B1(n2990), .B2(n36499), .ZN(
        n8994) );
  OAI22_X1 U2831 ( .A1(n38586), .A2(n38790), .B1(n2990), .B2(n36503), .ZN(
        n8995) );
  OAI22_X1 U2832 ( .A1(n38586), .A2(n38797), .B1(n2990), .B2(n36507), .ZN(
        n8996) );
  OAI22_X1 U2833 ( .A1(n38586), .A2(n38804), .B1(n2990), .B2(n36511), .ZN(
        n8997) );
  OAI22_X1 U2834 ( .A1(n38586), .A2(n38811), .B1(n2990), .B2(n36515), .ZN(
        n8998) );
  OAI22_X1 U2835 ( .A1(n38587), .A2(n38818), .B1(n2990), .B2(n36519), .ZN(
        n8999) );
  OAI22_X1 U2836 ( .A1(n38587), .A2(n38825), .B1(n38582), .B2(n36523), .ZN(
        n9000) );
  OAI22_X1 U2837 ( .A1(n38587), .A2(n38832), .B1(n38582), .B2(n36527), .ZN(
        n9001) );
  OAI22_X1 U2838 ( .A1(n38587), .A2(n38839), .B1(n38582), .B2(n36531), .ZN(
        n9002) );
  OAI22_X1 U2839 ( .A1(n38595), .A2(n38678), .B1(n38594), .B2(n35927), .ZN(
        n9011) );
  OAI22_X1 U2840 ( .A1(n38595), .A2(n38685), .B1(n38594), .B2(n35931), .ZN(
        n9012) );
  OAI22_X1 U2841 ( .A1(n38595), .A2(n38692), .B1(n38594), .B2(n35935), .ZN(
        n9013) );
  OAI22_X1 U2842 ( .A1(n38595), .A2(n38699), .B1(n38594), .B2(n35939), .ZN(
        n9014) );
  OAI22_X1 U2843 ( .A1(n38595), .A2(n38706), .B1(n38594), .B2(n35943), .ZN(
        n9015) );
  OAI22_X1 U2844 ( .A1(n38596), .A2(n38713), .B1(n38594), .B2(n35947), .ZN(
        n9016) );
  OAI22_X1 U2845 ( .A1(n38596), .A2(n38720), .B1(n38594), .B2(n35951), .ZN(
        n9017) );
  OAI22_X1 U2846 ( .A1(n38596), .A2(n38727), .B1(n38594), .B2(n35955), .ZN(
        n9018) );
  OAI22_X1 U2847 ( .A1(n38596), .A2(n38734), .B1(n38594), .B2(n35959), .ZN(
        n9019) );
  OAI22_X1 U2848 ( .A1(n38596), .A2(n38741), .B1(n38594), .B2(n35963), .ZN(
        n9020) );
  OAI22_X1 U2849 ( .A1(n38597), .A2(n38748), .B1(n38594), .B2(n35967), .ZN(
        n9021) );
  OAI22_X1 U2850 ( .A1(n38597), .A2(n38755), .B1(n38594), .B2(n35971), .ZN(
        n9022) );
  OAI22_X1 U2851 ( .A1(n38597), .A2(n38762), .B1(n38594), .B2(n35975), .ZN(
        n9023) );
  OAI22_X1 U2852 ( .A1(n38597), .A2(n38769), .B1(n38594), .B2(n35979), .ZN(
        n9024) );
  OAI22_X1 U2853 ( .A1(n38597), .A2(n38776), .B1(n2955), .B2(n35983), .ZN(
        n9025) );
  OAI22_X1 U2854 ( .A1(n38598), .A2(n38783), .B1(n2955), .B2(n35987), .ZN(
        n9026) );
  OAI22_X1 U2855 ( .A1(n38598), .A2(n38790), .B1(n2955), .B2(n35991), .ZN(
        n9027) );
  OAI22_X1 U2856 ( .A1(n38598), .A2(n38797), .B1(n2955), .B2(n35995), .ZN(
        n9028) );
  OAI22_X1 U2857 ( .A1(n38598), .A2(n38804), .B1(n2955), .B2(n35999), .ZN(
        n9029) );
  OAI22_X1 U2858 ( .A1(n38598), .A2(n38811), .B1(n2955), .B2(n36003), .ZN(
        n9030) );
  OAI22_X1 U2859 ( .A1(n38599), .A2(n38818), .B1(n2955), .B2(n36007), .ZN(
        n9031) );
  OAI22_X1 U2860 ( .A1(n38599), .A2(n38825), .B1(n38594), .B2(n36011), .ZN(
        n9032) );
  OAI22_X1 U2861 ( .A1(n38599), .A2(n38832), .B1(n38594), .B2(n36015), .ZN(
        n9033) );
  OAI22_X1 U2862 ( .A1(n38599), .A2(n38839), .B1(n38594), .B2(n36019), .ZN(
        n9034) );
  OAI22_X1 U2863 ( .A1(n38631), .A2(n38678), .B1(n38630), .B2(n35318), .ZN(
        n9107) );
  OAI22_X1 U2864 ( .A1(n38631), .A2(n38685), .B1(n38630), .B2(n35319), .ZN(
        n9108) );
  OAI22_X1 U2865 ( .A1(n38631), .A2(n38692), .B1(n38630), .B2(n35320), .ZN(
        n9109) );
  OAI22_X1 U2866 ( .A1(n38631), .A2(n38699), .B1(n38630), .B2(n35321), .ZN(
        n9110) );
  OAI22_X1 U2867 ( .A1(n38631), .A2(n38706), .B1(n38630), .B2(n35322), .ZN(
        n9111) );
  OAI22_X1 U2868 ( .A1(n38632), .A2(n38713), .B1(n38630), .B2(n35323), .ZN(
        n9112) );
  OAI22_X1 U2869 ( .A1(n38632), .A2(n38720), .B1(n38630), .B2(n35324), .ZN(
        n9113) );
  OAI22_X1 U2870 ( .A1(n38632), .A2(n38727), .B1(n38630), .B2(n35325), .ZN(
        n9114) );
  OAI22_X1 U2871 ( .A1(n38632), .A2(n38734), .B1(n38630), .B2(n35326), .ZN(
        n9115) );
  OAI22_X1 U2872 ( .A1(n38632), .A2(n38741), .B1(n38630), .B2(n35327), .ZN(
        n9116) );
  OAI22_X1 U2873 ( .A1(n38633), .A2(n38748), .B1(n38630), .B2(n35328), .ZN(
        n9117) );
  OAI22_X1 U2874 ( .A1(n38633), .A2(n38755), .B1(n38630), .B2(n35329), .ZN(
        n9118) );
  OAI22_X1 U2875 ( .A1(n38633), .A2(n38762), .B1(n38630), .B2(n35330), .ZN(
        n9119) );
  OAI22_X1 U2876 ( .A1(n38633), .A2(n38769), .B1(n38630), .B2(n35331), .ZN(
        n9120) );
  OAI22_X1 U2877 ( .A1(n38633), .A2(n38776), .B1(n2850), .B2(n35332), .ZN(
        n9121) );
  OAI22_X1 U2878 ( .A1(n38634), .A2(n38783), .B1(n2850), .B2(n35333), .ZN(
        n9122) );
  OAI22_X1 U2879 ( .A1(n38634), .A2(n38790), .B1(n2850), .B2(n35334), .ZN(
        n9123) );
  OAI22_X1 U2880 ( .A1(n38634), .A2(n38797), .B1(n2850), .B2(n35335), .ZN(
        n9124) );
  OAI22_X1 U2881 ( .A1(n38634), .A2(n38804), .B1(n2850), .B2(n35336), .ZN(
        n9125) );
  OAI22_X1 U2882 ( .A1(n38634), .A2(n38811), .B1(n2850), .B2(n35337), .ZN(
        n9126) );
  OAI22_X1 U2883 ( .A1(n38635), .A2(n38818), .B1(n2850), .B2(n35338), .ZN(
        n9127) );
  OAI22_X1 U2884 ( .A1(n38635), .A2(n38825), .B1(n38630), .B2(n35339), .ZN(
        n9128) );
  OAI22_X1 U2885 ( .A1(n38635), .A2(n38832), .B1(n38630), .B2(n35340), .ZN(
        n9129) );
  OAI22_X1 U2886 ( .A1(n38635), .A2(n38839), .B1(n38630), .B2(n35341), .ZN(
        n9130) );
  OAI22_X1 U2887 ( .A1(n38643), .A2(n38678), .B1(n38642), .B2(n36342), .ZN(
        n9139) );
  OAI22_X1 U2888 ( .A1(n38643), .A2(n38685), .B1(n38642), .B2(n36343), .ZN(
        n9140) );
  OAI22_X1 U2889 ( .A1(n38643), .A2(n38692), .B1(n38642), .B2(n36344), .ZN(
        n9141) );
  OAI22_X1 U2890 ( .A1(n38643), .A2(n38699), .B1(n38642), .B2(n36345), .ZN(
        n9142) );
  OAI22_X1 U2891 ( .A1(n38643), .A2(n38706), .B1(n38642), .B2(n36346), .ZN(
        n9143) );
  OAI22_X1 U2892 ( .A1(n38644), .A2(n38713), .B1(n38642), .B2(n36347), .ZN(
        n9144) );
  OAI22_X1 U2893 ( .A1(n38644), .A2(n38720), .B1(n38642), .B2(n36348), .ZN(
        n9145) );
  OAI22_X1 U2894 ( .A1(n38644), .A2(n38727), .B1(n38642), .B2(n36349), .ZN(
        n9146) );
  OAI22_X1 U2895 ( .A1(n38644), .A2(n38734), .B1(n38642), .B2(n36350), .ZN(
        n9147) );
  OAI22_X1 U2896 ( .A1(n38644), .A2(n38741), .B1(n38642), .B2(n36351), .ZN(
        n9148) );
  OAI22_X1 U2897 ( .A1(n38645), .A2(n38748), .B1(n38642), .B2(n36352), .ZN(
        n9149) );
  OAI22_X1 U2898 ( .A1(n38645), .A2(n38755), .B1(n38642), .B2(n36353), .ZN(
        n9150) );
  OAI22_X1 U2899 ( .A1(n38645), .A2(n38762), .B1(n2815), .B2(n36354), .ZN(
        n9151) );
  OAI22_X1 U2900 ( .A1(n38645), .A2(n38769), .B1(n2815), .B2(n36355), .ZN(
        n9152) );
  OAI22_X1 U2901 ( .A1(n38645), .A2(n38776), .B1(n2815), .B2(n36356), .ZN(
        n9153) );
  OAI22_X1 U2902 ( .A1(n38646), .A2(n38783), .B1(n2815), .B2(n36357), .ZN(
        n9154) );
  OAI22_X1 U2903 ( .A1(n38646), .A2(n38790), .B1(n2815), .B2(n36358), .ZN(
        n9155) );
  OAI22_X1 U2904 ( .A1(n38646), .A2(n38797), .B1(n2815), .B2(n36359), .ZN(
        n9156) );
  OAI22_X1 U2905 ( .A1(n38646), .A2(n38804), .B1(n2815), .B2(n36360), .ZN(
        n9157) );
  OAI22_X1 U2906 ( .A1(n38646), .A2(n38811), .B1(n2815), .B2(n36361), .ZN(
        n9158) );
  OAI22_X1 U2907 ( .A1(n38647), .A2(n38818), .B1(n2815), .B2(n36362), .ZN(
        n9159) );
  OAI22_X1 U2908 ( .A1(n38647), .A2(n38825), .B1(n38642), .B2(n36363), .ZN(
        n9160) );
  OAI22_X1 U2909 ( .A1(n38647), .A2(n38832), .B1(n38642), .B2(n36364), .ZN(
        n9161) );
  OAI22_X1 U2910 ( .A1(n38647), .A2(n38839), .B1(n38642), .B2(n36365), .ZN(
        n9162) );
  OAI22_X1 U2911 ( .A1(n38655), .A2(n38678), .B1(n38654), .B2(n35830), .ZN(
        n9171) );
  OAI22_X1 U2912 ( .A1(n38655), .A2(n38685), .B1(n38654), .B2(n35831), .ZN(
        n9172) );
  OAI22_X1 U2913 ( .A1(n38655), .A2(n38692), .B1(n38654), .B2(n35832), .ZN(
        n9173) );
  OAI22_X1 U2914 ( .A1(n38655), .A2(n38699), .B1(n38654), .B2(n35833), .ZN(
        n9174) );
  OAI22_X1 U2915 ( .A1(n38655), .A2(n38706), .B1(n38654), .B2(n35834), .ZN(
        n9175) );
  OAI22_X1 U2916 ( .A1(n38656), .A2(n38713), .B1(n38654), .B2(n35835), .ZN(
        n9176) );
  OAI22_X1 U2917 ( .A1(n38656), .A2(n38720), .B1(n38654), .B2(n35836), .ZN(
        n9177) );
  OAI22_X1 U2918 ( .A1(n38656), .A2(n38727), .B1(n38654), .B2(n35837), .ZN(
        n9178) );
  OAI22_X1 U2919 ( .A1(n38656), .A2(n38734), .B1(n38654), .B2(n35838), .ZN(
        n9179) );
  OAI22_X1 U2920 ( .A1(n38656), .A2(n38741), .B1(n38654), .B2(n35839), .ZN(
        n9180) );
  OAI22_X1 U2921 ( .A1(n38657), .A2(n38748), .B1(n38654), .B2(n35840), .ZN(
        n9181) );
  OAI22_X1 U2922 ( .A1(n38657), .A2(n38755), .B1(n38654), .B2(n35841), .ZN(
        n9182) );
  OAI22_X1 U2923 ( .A1(n38657), .A2(n38762), .B1(n2778), .B2(n35842), .ZN(
        n9183) );
  OAI22_X1 U2924 ( .A1(n38657), .A2(n38769), .B1(n2778), .B2(n35843), .ZN(
        n9184) );
  OAI22_X1 U2925 ( .A1(n38657), .A2(n38776), .B1(n2778), .B2(n35844), .ZN(
        n9185) );
  OAI22_X1 U2926 ( .A1(n38658), .A2(n38783), .B1(n2778), .B2(n35845), .ZN(
        n9186) );
  OAI22_X1 U2927 ( .A1(n38658), .A2(n38790), .B1(n2778), .B2(n35846), .ZN(
        n9187) );
  OAI22_X1 U2928 ( .A1(n38658), .A2(n38797), .B1(n2778), .B2(n35847), .ZN(
        n9188) );
  OAI22_X1 U2929 ( .A1(n38658), .A2(n38804), .B1(n2778), .B2(n35848), .ZN(
        n9189) );
  OAI22_X1 U2930 ( .A1(n38658), .A2(n38811), .B1(n2778), .B2(n35849), .ZN(
        n9190) );
  OAI22_X1 U2931 ( .A1(n38659), .A2(n38818), .B1(n2778), .B2(n35850), .ZN(
        n9191) );
  OAI22_X1 U2932 ( .A1(n38659), .A2(n38825), .B1(n38654), .B2(n35851), .ZN(
        n9192) );
  OAI22_X1 U2933 ( .A1(n38659), .A2(n38832), .B1(n38654), .B2(n35852), .ZN(
        n9193) );
  OAI22_X1 U2934 ( .A1(n38659), .A2(n38839), .B1(n38654), .B2(n35853), .ZN(
        n9194) );
  BUF_X1 U2935 ( .A(n38914), .Z(n38913) );
  BUF_X1 U2936 ( .A(n38915), .Z(n38911) );
  BUF_X1 U2937 ( .A(n38915), .Z(n38912) );
  BUF_X1 U2938 ( .A(n3303), .Z(n38480) );
  BUF_X1 U2939 ( .A(n3303), .Z(n38481) );
  INV_X1 U2940 ( .A(n2778), .ZN(n38662) );
  OAI21_X1 U2941 ( .B1(n38653), .B2(n2812), .A(n38919), .ZN(n2778) );
  INV_X1 U2942 ( .A(n3200), .ZN(n38518) );
  OAI21_X1 U2943 ( .B1(n2812), .B2(n38507), .A(n38917), .ZN(n3200) );
  INV_X1 U2944 ( .A(n3165), .ZN(n38530) );
  OAI21_X1 U2945 ( .B1(n2812), .B2(n38521), .A(n38917), .ZN(n3165) );
  INV_X1 U2946 ( .A(n3130), .ZN(n38542) );
  OAI21_X1 U2947 ( .B1(n2812), .B2(n38531), .A(n38917), .ZN(n3130) );
  INV_X1 U2948 ( .A(n3025), .ZN(n38578) );
  OAI21_X1 U2949 ( .B1(n2812), .B2(n38567), .A(n38917), .ZN(n3025) );
  INV_X1 U2950 ( .A(n2990), .ZN(n38590) );
  OAI21_X1 U2951 ( .B1(n2812), .B2(n38581), .A(n38917), .ZN(n2990) );
  INV_X1 U2952 ( .A(n2955), .ZN(n38602) );
  OAI21_X1 U2953 ( .B1(n2812), .B2(n38591), .A(n38920), .ZN(n2955) );
  INV_X1 U2954 ( .A(n2850), .ZN(n38638) );
  OAI21_X1 U2955 ( .B1(n2812), .B2(n38627), .A(n38919), .ZN(n2850) );
  INV_X1 U2956 ( .A(n2815), .ZN(n38650) );
  OAI21_X1 U2957 ( .B1(n2812), .B2(n38641), .A(n38917), .ZN(n2815) );
  INV_X1 U2958 ( .A(n5474), .ZN(n37813) );
  OAI21_X1 U2959 ( .B1(n5016), .B2(n5507), .A(n38917), .ZN(n5474) );
  INV_X1 U2960 ( .A(n5439), .ZN(n37825) );
  OAI21_X1 U2961 ( .B1(n5016), .B2(n37814), .A(n38917), .ZN(n5439) );
  INV_X1 U2962 ( .A(n5404), .ZN(n37837) );
  OAI21_X1 U2963 ( .B1(n5016), .B2(n37828), .A(n38920), .ZN(n5404) );
  INV_X1 U2964 ( .A(n5369), .ZN(n37849) );
  OAI21_X1 U2965 ( .B1(n5016), .B2(n37838), .A(n38917), .ZN(n5369) );
  INV_X1 U2966 ( .A(n5334), .ZN(n37858) );
  OAI21_X1 U2967 ( .B1(n5016), .B2(n5367), .A(n38916), .ZN(n5334) );
  INV_X1 U2968 ( .A(n5299), .ZN(n37867) );
  OAI21_X1 U2969 ( .B1(n5016), .B2(n5332), .A(n38917), .ZN(n5299) );
  INV_X1 U2970 ( .A(n5264), .ZN(n37879) );
  OAI21_X1 U2971 ( .B1(n5016), .B2(n37868), .A(n38919), .ZN(n5264) );
  INV_X1 U2972 ( .A(n5229), .ZN(n37891) );
  OAI21_X1 U2973 ( .B1(n5016), .B2(n37882), .A(n38920), .ZN(n5229) );
  INV_X1 U2974 ( .A(n5194), .ZN(n37903) );
  OAI21_X1 U2975 ( .B1(n5016), .B2(n37892), .A(n38920), .ZN(n5194) );
  INV_X1 U2976 ( .A(n5159), .ZN(n37912) );
  OAI21_X1 U2977 ( .B1(n5016), .B2(n5192), .A(n38919), .ZN(n5159) );
  INV_X1 U2978 ( .A(n5124), .ZN(n37921) );
  OAI21_X1 U2979 ( .B1(n5016), .B2(n5157), .A(n38918), .ZN(n5124) );
  INV_X1 U2980 ( .A(n5089), .ZN(n37933) );
  OAI21_X1 U2981 ( .B1(n5016), .B2(n37922), .A(n38918), .ZN(n5089) );
  INV_X1 U2982 ( .A(n5054), .ZN(n37945) );
  OAI21_X1 U2983 ( .B1(n5016), .B2(n37936), .A(n38918), .ZN(n5054) );
  INV_X1 U2984 ( .A(n5019), .ZN(n37957) );
  OAI21_X1 U2985 ( .B1(n5016), .B2(n37946), .A(n38919), .ZN(n5019) );
  INV_X1 U2986 ( .A(n4983), .ZN(n37966) );
  OAI21_X1 U2987 ( .B1(n5016), .B2(n5017), .A(n38920), .ZN(n4983) );
  NOR2_X2 U2988 ( .A1(n9630), .A2(n9629), .ZN(n9583) );
  BUF_X1 U2989 ( .A(n5437), .Z(n37828) );
  BUF_X1 U2990 ( .A(n5262), .Z(n37882) );
  BUF_X1 U2991 ( .A(n5087), .Z(n37936) );
  BUF_X1 U2992 ( .A(n5472), .Z(n37816) );
  BUF_X1 U2993 ( .A(n5297), .Z(n37870) );
  BUF_X1 U2994 ( .A(n5122), .Z(n37924) );
  BUF_X1 U2995 ( .A(n5437), .Z(n37826) );
  BUF_X1 U2996 ( .A(n5262), .Z(n37880) );
  BUF_X1 U2997 ( .A(n5087), .Z(n37934) );
  BUF_X1 U2998 ( .A(n5437), .Z(n37827) );
  BUF_X1 U2999 ( .A(n5262), .Z(n37881) );
  BUF_X1 U3000 ( .A(n5087), .Z(n37935) );
  BUF_X1 U3001 ( .A(n5402), .Z(n37840) );
  BUF_X1 U3002 ( .A(n5227), .Z(n37894) );
  BUF_X1 U3003 ( .A(n5052), .Z(n37948) );
  BUF_X1 U3004 ( .A(n5472), .Z(n37814) );
  BUF_X1 U3005 ( .A(n5297), .Z(n37868) );
  BUF_X1 U3006 ( .A(n5122), .Z(n37922) );
  BUF_X1 U3007 ( .A(n5472), .Z(n37815) );
  BUF_X1 U3008 ( .A(n5297), .Z(n37869) );
  BUF_X1 U3009 ( .A(n5122), .Z(n37923) );
  BUF_X1 U3010 ( .A(n5402), .Z(n37838) );
  BUF_X1 U3011 ( .A(n5227), .Z(n37892) );
  BUF_X1 U3012 ( .A(n5052), .Z(n37946) );
  BUF_X1 U3013 ( .A(n5402), .Z(n37839) );
  BUF_X1 U3014 ( .A(n5227), .Z(n37893) );
  BUF_X1 U3015 ( .A(n5052), .Z(n37947) );
  AND3_X1 U3016 ( .A1(n9604), .A2(n9603), .A3(n9625), .ZN(n9581) );
  AND3_X1 U3017 ( .A1(n9604), .A2(n9614), .A3(n9619), .ZN(n9578) );
  AND3_X1 U3018 ( .A1(n9604), .A2(n9603), .A3(n9601), .ZN(n9589) );
  AND3_X1 U3019 ( .A1(n9604), .A2(n9614), .A3(n9615), .ZN(n9574) );
  NAND2_X1 U3020 ( .A1(n9585), .A2(n9584), .ZN(n3934) );
  NAND2_X1 U3021 ( .A1(n9586), .A2(n9587), .ZN(n3339) );
  NAND2_X1 U3022 ( .A1(n9585), .A2(n9589), .ZN(n3864) );
  NAND2_X1 U3023 ( .A1(n9586), .A2(n9589), .ZN(n3304) );
  NAND2_X1 U3024 ( .A1(n9585), .A2(n9571), .ZN(n4316) );
  NAND2_X1 U3025 ( .A1(n9586), .A2(n9573), .ZN(n3689) );
  NAND2_X1 U3026 ( .A1(n9585), .A2(n9574), .ZN(n4246) );
  NAND2_X1 U3027 ( .A1(n9586), .A2(n9574), .ZN(n3654) );
  NAND2_X1 U3028 ( .A1(n9585), .A2(n9590), .ZN(n4421) );
  NAND2_X1 U3029 ( .A1(n9586), .A2(n9590), .ZN(n3829) );
  NAND2_X1 U3030 ( .A1(n9586), .A2(n9572), .ZN(n3759) );
  NAND2_X1 U3031 ( .A1(n9585), .A2(n9572), .ZN(n4351) );
  NAND2_X1 U3032 ( .A1(n9585), .A2(n9580), .ZN(n4039) );
  NAND2_X1 U3033 ( .A1(n9586), .A2(n9580), .ZN(n3479) );
  NAND2_X1 U3034 ( .A1(n9586), .A2(n9599), .ZN(n3409) );
  NAND2_X1 U3035 ( .A1(n9585), .A2(n9599), .ZN(n3969) );
  NAND2_X1 U3036 ( .A1(n9586), .A2(n9578), .ZN(n3584) );
  NAND2_X1 U3037 ( .A1(n9585), .A2(n9578), .ZN(n4176) );
  NAND2_X1 U3038 ( .A1(n9585), .A2(n9577), .ZN(n4136) );
  NAND2_X1 U3039 ( .A1(n9586), .A2(n9579), .ZN(n3514) );
  NAND2_X1 U3040 ( .A1(n9583), .A2(n9584), .ZN(n4526) );
  NAND2_X1 U3041 ( .A1(n9583), .A2(n9571), .ZN(n4876) );
  NAND2_X1 U3042 ( .A1(n9583), .A2(n9590), .ZN(n4981) );
  NAND2_X1 U3043 ( .A1(n9583), .A2(n9591), .ZN(n4946) );
  NAND2_X1 U3044 ( .A1(n9583), .A2(n9580), .ZN(n4631) );
  NAND2_X1 U3045 ( .A1(n9583), .A2(n9575), .ZN(n4771) );
  NAND2_X1 U3046 ( .A1(n9583), .A2(n9577), .ZN(n4701) );
  NAND2_X1 U3047 ( .A1(n9578), .A2(n9597), .ZN(n3023) );
  NAND2_X1 U3048 ( .A1(n9575), .A2(n9597), .ZN(n3058) );
  NAND2_X1 U3049 ( .A1(n9577), .A2(n9597), .ZN(n2988) );
  NAND2_X1 U3050 ( .A1(n9599), .A2(n9597), .ZN(n2848) );
  NAND2_X1 U3051 ( .A1(n9581), .A2(n9597), .ZN(n2883) );
  NAND2_X1 U3052 ( .A1(n9584), .A2(n9597), .ZN(n2811) );
  NAND2_X1 U3053 ( .A1(n9572), .A2(n9597), .ZN(n3198) );
  NAND2_X1 U3054 ( .A1(n9591), .A2(n9597), .ZN(n3233) );
  NAND2_X1 U3055 ( .A1(n9571), .A2(n9597), .ZN(n3163) );
  NAND2_X1 U3056 ( .A1(n9585), .A2(n9587), .ZN(n3899) );
  NAND2_X1 U3057 ( .A1(n9585), .A2(n9573), .ZN(n4281) );
  NAND2_X1 U3058 ( .A1(n9586), .A2(n9575), .ZN(n3619) );
  NAND2_X1 U3059 ( .A1(n9585), .A2(n9575), .ZN(n4211) );
  NAND2_X1 U3060 ( .A1(n9586), .A2(n9591), .ZN(n3794) );
  NAND2_X1 U3061 ( .A1(n9585), .A2(n9591), .ZN(n4386) );
  NAND2_X1 U3062 ( .A1(n9586), .A2(n9571), .ZN(n3724) );
  NAND2_X1 U3063 ( .A1(n9586), .A2(n9581), .ZN(n3444) );
  NAND2_X1 U3064 ( .A1(n9585), .A2(n9581), .ZN(n4004) );
  NAND2_X1 U3065 ( .A1(n9586), .A2(n9584), .ZN(n3374) );
  NAND2_X1 U3066 ( .A1(n9586), .A2(n9577), .ZN(n3549) );
  NAND2_X1 U3067 ( .A1(n9585), .A2(n9579), .ZN(n4074) );
  NAND2_X1 U3068 ( .A1(n9583), .A2(n9587), .ZN(n4491) );
  NAND2_X1 U3069 ( .A1(n9583), .A2(n9573), .ZN(n4841) );
  NAND2_X1 U3070 ( .A1(n9583), .A2(n9572), .ZN(n4911) );
  NAND2_X1 U3071 ( .A1(n9583), .A2(n9599), .ZN(n4561) );
  NAND2_X1 U3072 ( .A1(n9583), .A2(n9579), .ZN(n4666) );
  AND2_X1 U3073 ( .A1(n9590), .A2(n9597), .ZN(n3268) );
  AND2_X1 U3074 ( .A1(n9573), .A2(n9597), .ZN(n3128) );
  AND2_X1 U3075 ( .A1(n9574), .A2(n9597), .ZN(n3093) );
  AND2_X1 U3076 ( .A1(n9579), .A2(n9597), .ZN(n2953) );
  AND2_X1 U3077 ( .A1(n9580), .A2(n9597), .ZN(n2918) );
  AND2_X1 U3078 ( .A1(n9587), .A2(n9597), .ZN(n2776) );
  AND2_X1 U3079 ( .A1(n9589), .A2(n9597), .ZN(n2740) );
  INV_X1 U3080 ( .A(n5157), .ZN(n5525) );
  INV_X1 U3081 ( .A(n5332), .ZN(n5522) );
  INV_X1 U3082 ( .A(n5507), .ZN(n5531) );
  INV_X1 U3083 ( .A(n5367), .ZN(n5523) );
  INV_X1 U3084 ( .A(n5192), .ZN(n5526) );
  INV_X1 U3085 ( .A(n5017), .ZN(n5540) );
  INV_X1 U3086 ( .A(n9560), .ZN(n5532) );
  NAND2_X1 U3087 ( .A1(WR_enable), .A2(ENABLE), .ZN(n2812) );
  AOI221_X1 U3088 ( .B1(net253671), .B2(n37784), .C1(net253639), .C2(n37781), 
        .A(n5841), .ZN(n5840) );
  OAI222_X1 U3089 ( .A1(n37838), .A2(n35854), .B1(n37814), .B2(n35342), .C1(
        n37828), .C2(n36366), .ZN(n5841) );
  AOI221_X1 U3090 ( .B1(net253799), .B2(n37757), .C1(net253991), .C2(n37754), 
        .A(n5859), .ZN(n5857) );
  OAI222_X1 U3091 ( .A1(n38357), .A2(n35855), .B1(n38174), .B2(n35343), .C1(
        n38002), .C2(n36367), .ZN(n5859) );
  AOI221_X1 U3092 ( .B1(net254023), .B2(n37751), .C1(net254215), .C2(n37748), 
        .A(n5861), .ZN(n5855) );
  OAI222_X1 U3093 ( .A1(n38021), .A2(n35856), .B1(n38369), .B2(n35344), .C1(
        n38197), .C2(n36368), .ZN(n5861) );
  AOI221_X1 U3094 ( .B1(net253959), .B2(n37745), .C1(net254151), .C2(n37742), 
        .A(n5863), .ZN(n5854) );
  OAI222_X1 U3095 ( .A1(n37967), .A2(n35857), .B1(n38315), .B2(n35345), .C1(
        n38143), .C2(n36369), .ZN(n5863) );
  AOI221_X1 U3096 ( .B1(net254183), .B2(n37739), .C1(net253767), .C2(n37736), 
        .A(n5864), .ZN(n5853) );
  OAI222_X1 U3097 ( .A1(n38162), .A2(n35858), .B1(n37979), .B2(n35346), .C1(
        n38338), .C2(n36370), .ZN(n5864) );
  AOI221_X1 U3098 ( .B1(net254087), .B2(n37733), .C1(net254279), .C2(n37730), 
        .A(n5869), .ZN(n5868) );
  OAI222_X1 U3099 ( .A1(n38075), .A2(n35859), .B1(n38423), .B2(n35347), .C1(
        n38251), .C2(n36371), .ZN(n5869) );
  AOI221_X1 U3100 ( .B1(net254311), .B2(n37727), .C1(net253895), .C2(n37724), 
        .A(n5870), .ZN(n5867) );
  OAI222_X1 U3101 ( .A1(n38270), .A2(n35860), .B1(n38087), .B2(n35348), .C1(
        n38446), .C2(n36372), .ZN(n5870) );
  AOI221_X1 U3102 ( .B1(net254247), .B2(n37721), .C1(net253831), .C2(n37718), 
        .A(n5871), .ZN(n5866) );
  OAI222_X1 U3103 ( .A1(n38216), .A2(n35861), .B1(n38033), .B2(n35349), .C1(
        n38392), .C2(n36373), .ZN(n5871) );
  AOI221_X1 U3104 ( .B1(net253863), .B2(n37715), .C1(net254055), .C2(n37712), 
        .A(n5872), .ZN(n5865) );
  OAI222_X1 U3105 ( .A1(n38411), .A2(n35862), .B1(n38228), .B2(n35350), .C1(
        n38056), .C2(n36374), .ZN(n5872) );
  AOI221_X1 U3106 ( .B1(net253672), .B2(n37784), .C1(net253640), .C2(n37781), 
        .A(n5799), .ZN(n5798) );
  OAI222_X1 U3107 ( .A1(n37838), .A2(n35863), .B1(n37814), .B2(n35351), .C1(
        n37828), .C2(n36375), .ZN(n5799) );
  AOI221_X1 U3108 ( .B1(net253800), .B2(n37757), .C1(net253992), .C2(n37754), 
        .A(n5817), .ZN(n5815) );
  OAI222_X1 U3109 ( .A1(n38357), .A2(n35864), .B1(n38174), .B2(n35352), .C1(
        n38002), .C2(n36376), .ZN(n5817) );
  AOI221_X1 U3110 ( .B1(net254024), .B2(n37751), .C1(net254216), .C2(n37748), 
        .A(n5819), .ZN(n5813) );
  OAI222_X1 U3111 ( .A1(n38021), .A2(n35865), .B1(n38369), .B2(n35353), .C1(
        n38197), .C2(n36377), .ZN(n5819) );
  AOI221_X1 U3112 ( .B1(net253960), .B2(n37745), .C1(net254152), .C2(n37742), 
        .A(n5821), .ZN(n5812) );
  OAI222_X1 U3113 ( .A1(n37967), .A2(n35866), .B1(n38315), .B2(n35354), .C1(
        n38143), .C2(n36378), .ZN(n5821) );
  AOI221_X1 U3114 ( .B1(net254184), .B2(n37739), .C1(net253768), .C2(n37736), 
        .A(n5822), .ZN(n5811) );
  OAI222_X1 U3115 ( .A1(n38162), .A2(n35867), .B1(n37979), .B2(n35355), .C1(
        n38338), .C2(n36379), .ZN(n5822) );
  AOI221_X1 U3116 ( .B1(net254088), .B2(n37733), .C1(net254280), .C2(n37730), 
        .A(n5827), .ZN(n5826) );
  OAI222_X1 U3117 ( .A1(n38075), .A2(n35868), .B1(n38423), .B2(n35356), .C1(
        n38251), .C2(n36380), .ZN(n5827) );
  AOI221_X1 U3118 ( .B1(net254312), .B2(n37727), .C1(net253896), .C2(n37724), 
        .A(n5828), .ZN(n5825) );
  OAI222_X1 U3119 ( .A1(n38270), .A2(n35869), .B1(n38087), .B2(n35357), .C1(
        n38446), .C2(n36381), .ZN(n5828) );
  AOI221_X1 U3120 ( .B1(net254248), .B2(n37721), .C1(net253832), .C2(n37718), 
        .A(n5829), .ZN(n5824) );
  OAI222_X1 U3121 ( .A1(n38216), .A2(n35870), .B1(n38033), .B2(n35358), .C1(
        n38392), .C2(n36382), .ZN(n5829) );
  AOI221_X1 U3122 ( .B1(net253864), .B2(n37715), .C1(net254056), .C2(n37712), 
        .A(n5830), .ZN(n5823) );
  OAI222_X1 U3123 ( .A1(n38411), .A2(n35871), .B1(n38228), .B2(n35359), .C1(
        n38056), .C2(n36383), .ZN(n5830) );
  AOI221_X1 U3124 ( .B1(net253673), .B2(n37784), .C1(net253641), .C2(n37781), 
        .A(n5757), .ZN(n5756) );
  OAI222_X1 U3125 ( .A1(n37838), .A2(n35872), .B1(n37814), .B2(n35360), .C1(
        n37828), .C2(n36384), .ZN(n5757) );
  AOI221_X1 U3126 ( .B1(net253801), .B2(n37757), .C1(net253993), .C2(n37754), 
        .A(n5775), .ZN(n5773) );
  OAI222_X1 U3127 ( .A1(n38357), .A2(n35873), .B1(n38174), .B2(n35361), .C1(
        n38002), .C2(n36385), .ZN(n5775) );
  AOI221_X1 U3128 ( .B1(net254025), .B2(n37751), .C1(net254217), .C2(n37748), 
        .A(n5777), .ZN(n5771) );
  OAI222_X1 U3129 ( .A1(n38021), .A2(n35874), .B1(n38369), .B2(n35362), .C1(
        n38197), .C2(n36386), .ZN(n5777) );
  AOI221_X1 U3130 ( .B1(net253961), .B2(n37745), .C1(net254153), .C2(n37742), 
        .A(n5779), .ZN(n5770) );
  OAI222_X1 U3131 ( .A1(n37967), .A2(n35875), .B1(n38315), .B2(n35363), .C1(
        n38143), .C2(n36387), .ZN(n5779) );
  AOI221_X1 U3132 ( .B1(net254185), .B2(n37739), .C1(net253769), .C2(n37736), 
        .A(n5780), .ZN(n5769) );
  OAI222_X1 U3133 ( .A1(n38162), .A2(n35876), .B1(n37979), .B2(n35364), .C1(
        n38338), .C2(n36388), .ZN(n5780) );
  AOI221_X1 U3134 ( .B1(net254089), .B2(n37733), .C1(net254281), .C2(n37730), 
        .A(n5785), .ZN(n5784) );
  OAI222_X1 U3135 ( .A1(n38075), .A2(n35877), .B1(n38423), .B2(n35365), .C1(
        n38251), .C2(n36389), .ZN(n5785) );
  AOI221_X1 U3136 ( .B1(net254313), .B2(n37727), .C1(net253897), .C2(n37724), 
        .A(n5786), .ZN(n5783) );
  OAI222_X1 U3137 ( .A1(n38270), .A2(n35878), .B1(n38087), .B2(n35366), .C1(
        n38446), .C2(n36390), .ZN(n5786) );
  AOI221_X1 U3138 ( .B1(net254249), .B2(n37721), .C1(net253833), .C2(n37718), 
        .A(n5787), .ZN(n5782) );
  OAI222_X1 U3139 ( .A1(n38216), .A2(n35879), .B1(n38033), .B2(n35367), .C1(
        n38392), .C2(n36391), .ZN(n5787) );
  AOI221_X1 U3140 ( .B1(net253865), .B2(n37715), .C1(net254057), .C2(n37712), 
        .A(n5788), .ZN(n5781) );
  OAI222_X1 U3141 ( .A1(n38411), .A2(n35880), .B1(n38228), .B2(n35368), .C1(
        n38056), .C2(n36392), .ZN(n5788) );
  AOI221_X1 U3142 ( .B1(net253674), .B2(n37784), .C1(net253642), .C2(n37781), 
        .A(n5715), .ZN(n5714) );
  OAI222_X1 U3143 ( .A1(n37838), .A2(n35881), .B1(n37814), .B2(n35369), .C1(
        n37828), .C2(n36393), .ZN(n5715) );
  AOI221_X1 U3144 ( .B1(net253802), .B2(n37757), .C1(net253994), .C2(n37754), 
        .A(n5733), .ZN(n5731) );
  OAI222_X1 U3145 ( .A1(n38357), .A2(n35882), .B1(n38174), .B2(n35370), .C1(
        n38002), .C2(n36394), .ZN(n5733) );
  AOI221_X1 U3146 ( .B1(net254026), .B2(n37751), .C1(net254218), .C2(n37748), 
        .A(n5735), .ZN(n5729) );
  OAI222_X1 U3147 ( .A1(n38021), .A2(n35883), .B1(n38369), .B2(n35371), .C1(
        n38197), .C2(n36395), .ZN(n5735) );
  AOI221_X1 U3148 ( .B1(net253962), .B2(n37745), .C1(net254154), .C2(n37742), 
        .A(n5737), .ZN(n5728) );
  OAI222_X1 U3149 ( .A1(n37967), .A2(n35884), .B1(n38315), .B2(n35372), .C1(
        n38143), .C2(n36396), .ZN(n5737) );
  AOI221_X1 U3150 ( .B1(net254186), .B2(n37739), .C1(net253770), .C2(n37736), 
        .A(n5738), .ZN(n5727) );
  OAI222_X1 U3151 ( .A1(n38162), .A2(n35885), .B1(n37979), .B2(n35373), .C1(
        n38338), .C2(n36397), .ZN(n5738) );
  AOI221_X1 U3152 ( .B1(net254090), .B2(n37733), .C1(net254282), .C2(n37730), 
        .A(n5743), .ZN(n5742) );
  OAI222_X1 U3153 ( .A1(n38075), .A2(n35886), .B1(n38423), .B2(n35374), .C1(
        n38251), .C2(n36398), .ZN(n5743) );
  AOI221_X1 U3154 ( .B1(net254314), .B2(n37727), .C1(net253898), .C2(n37724), 
        .A(n5744), .ZN(n5741) );
  OAI222_X1 U3155 ( .A1(n38270), .A2(n35887), .B1(n38087), .B2(n35375), .C1(
        n38446), .C2(n36399), .ZN(n5744) );
  AOI221_X1 U3156 ( .B1(net254250), .B2(n37721), .C1(net253834), .C2(n37718), 
        .A(n5745), .ZN(n5740) );
  OAI222_X1 U3157 ( .A1(n38216), .A2(n35888), .B1(n38033), .B2(n35376), .C1(
        n38392), .C2(n36400), .ZN(n5745) );
  AOI221_X1 U3158 ( .B1(net253866), .B2(n37715), .C1(net254058), .C2(n37712), 
        .A(n5746), .ZN(n5739) );
  OAI222_X1 U3159 ( .A1(n38411), .A2(n35889), .B1(n38228), .B2(n35377), .C1(
        n38056), .C2(n36401), .ZN(n5746) );
  AOI221_X1 U3160 ( .B1(net253675), .B2(n37784), .C1(net253643), .C2(n37781), 
        .A(n5673), .ZN(n5672) );
  OAI222_X1 U3161 ( .A1(n37838), .A2(n35890), .B1(n37814), .B2(n35378), .C1(
        n37828), .C2(n36402), .ZN(n5673) );
  AOI221_X1 U3162 ( .B1(net253803), .B2(n37757), .C1(net253995), .C2(n37754), 
        .A(n5691), .ZN(n5689) );
  OAI222_X1 U3163 ( .A1(n38357), .A2(n35891), .B1(n38174), .B2(n35379), .C1(
        n38002), .C2(n36403), .ZN(n5691) );
  AOI221_X1 U3164 ( .B1(net254027), .B2(n37751), .C1(net254219), .C2(n37748), 
        .A(n5693), .ZN(n5687) );
  OAI222_X1 U3165 ( .A1(n38021), .A2(n35892), .B1(n38369), .B2(n35380), .C1(
        n38197), .C2(n36404), .ZN(n5693) );
  AOI221_X1 U3166 ( .B1(net253963), .B2(n37745), .C1(net254155), .C2(n37742), 
        .A(n5695), .ZN(n5686) );
  OAI222_X1 U3167 ( .A1(n37967), .A2(n35893), .B1(n38315), .B2(n35381), .C1(
        n38143), .C2(n36405), .ZN(n5695) );
  AOI221_X1 U3168 ( .B1(net254187), .B2(n37739), .C1(net253771), .C2(n37736), 
        .A(n5696), .ZN(n5685) );
  OAI222_X1 U3169 ( .A1(n38162), .A2(n35894), .B1(n37979), .B2(n35382), .C1(
        n38338), .C2(n36406), .ZN(n5696) );
  AOI221_X1 U3170 ( .B1(net254091), .B2(n37733), .C1(net254283), .C2(n37730), 
        .A(n5701), .ZN(n5700) );
  OAI222_X1 U3171 ( .A1(n38075), .A2(n35895), .B1(n38423), .B2(n35383), .C1(
        n38251), .C2(n36407), .ZN(n5701) );
  AOI221_X1 U3172 ( .B1(net254315), .B2(n37727), .C1(net253899), .C2(n37724), 
        .A(n5702), .ZN(n5699) );
  OAI222_X1 U3173 ( .A1(n38270), .A2(n35896), .B1(n38087), .B2(n35384), .C1(
        n38446), .C2(n36408), .ZN(n5702) );
  AOI221_X1 U3174 ( .B1(net254251), .B2(n37721), .C1(net253835), .C2(n37718), 
        .A(n5703), .ZN(n5698) );
  OAI222_X1 U3175 ( .A1(n38216), .A2(n35897), .B1(n38033), .B2(n35385), .C1(
        n38392), .C2(n36409), .ZN(n5703) );
  AOI221_X1 U3176 ( .B1(net253867), .B2(n37715), .C1(net254059), .C2(n37712), 
        .A(n5704), .ZN(n5697) );
  OAI222_X1 U3177 ( .A1(n38411), .A2(n35898), .B1(n38228), .B2(n35386), .C1(
        n38056), .C2(n36410), .ZN(n5704) );
  AOI221_X1 U3178 ( .B1(net253676), .B2(n37784), .C1(net253644), .C2(n37781), 
        .A(n5631), .ZN(n5630) );
  OAI222_X1 U3179 ( .A1(n37838), .A2(n35899), .B1(n37814), .B2(n35387), .C1(
        n37828), .C2(n36411), .ZN(n5631) );
  AOI221_X1 U3180 ( .B1(net253804), .B2(n37757), .C1(net253996), .C2(n37754), 
        .A(n5649), .ZN(n5647) );
  OAI222_X1 U3181 ( .A1(n38357), .A2(n35900), .B1(n38174), .B2(n35388), .C1(
        n38002), .C2(n36412), .ZN(n5649) );
  AOI221_X1 U3182 ( .B1(net254028), .B2(n37751), .C1(net254220), .C2(n37748), 
        .A(n5651), .ZN(n5645) );
  OAI222_X1 U3183 ( .A1(n38021), .A2(n35901), .B1(n38369), .B2(n35389), .C1(
        n38197), .C2(n36413), .ZN(n5651) );
  AOI221_X1 U3184 ( .B1(net253964), .B2(n37745), .C1(net254156), .C2(n37742), 
        .A(n5653), .ZN(n5644) );
  OAI222_X1 U3185 ( .A1(n37967), .A2(n35902), .B1(n38315), .B2(n35390), .C1(
        n38143), .C2(n36414), .ZN(n5653) );
  AOI221_X1 U3186 ( .B1(net254188), .B2(n37739), .C1(net253772), .C2(n37736), 
        .A(n5654), .ZN(n5643) );
  OAI222_X1 U3187 ( .A1(n38162), .A2(n35903), .B1(n37979), .B2(n35391), .C1(
        n38338), .C2(n36415), .ZN(n5654) );
  AOI221_X1 U3188 ( .B1(net254092), .B2(n37733), .C1(net254284), .C2(n37730), 
        .A(n5659), .ZN(n5658) );
  OAI222_X1 U3189 ( .A1(n38075), .A2(n35904), .B1(n38423), .B2(n35392), .C1(
        n38251), .C2(n36416), .ZN(n5659) );
  AOI221_X1 U3190 ( .B1(net254316), .B2(n37727), .C1(net253900), .C2(n37724), 
        .A(n5660), .ZN(n5657) );
  OAI222_X1 U3191 ( .A1(n38270), .A2(n35905), .B1(n38087), .B2(n35393), .C1(
        n38446), .C2(n36417), .ZN(n5660) );
  AOI221_X1 U3192 ( .B1(net254252), .B2(n37721), .C1(net253836), .C2(n37718), 
        .A(n5661), .ZN(n5656) );
  OAI222_X1 U3193 ( .A1(n38216), .A2(n35906), .B1(n38033), .B2(n35394), .C1(
        n38392), .C2(n36418), .ZN(n5661) );
  AOI221_X1 U3194 ( .B1(net253868), .B2(n37715), .C1(net254060), .C2(n37712), 
        .A(n5662), .ZN(n5655) );
  OAI222_X1 U3195 ( .A1(n38411), .A2(n35907), .B1(n38228), .B2(n35395), .C1(
        n38056), .C2(n36419), .ZN(n5662) );
  AOI221_X1 U3196 ( .B1(net253677), .B2(n37784), .C1(net253645), .C2(n37781), 
        .A(n5589), .ZN(n5588) );
  OAI222_X1 U3197 ( .A1(n37838), .A2(n35908), .B1(n37814), .B2(n35396), .C1(
        n37828), .C2(n36420), .ZN(n5589) );
  AOI221_X1 U3198 ( .B1(net253805), .B2(n37757), .C1(net253997), .C2(n37754), 
        .A(n5607), .ZN(n5605) );
  OAI222_X1 U3199 ( .A1(n38357), .A2(n35909), .B1(n38174), .B2(n35397), .C1(
        n38002), .C2(n36421), .ZN(n5607) );
  AOI221_X1 U3200 ( .B1(net254029), .B2(n37751), .C1(net254221), .C2(n37748), 
        .A(n5609), .ZN(n5603) );
  OAI222_X1 U3201 ( .A1(n38021), .A2(n35910), .B1(n38369), .B2(n35398), .C1(
        n38197), .C2(n36422), .ZN(n5609) );
  AOI221_X1 U3202 ( .B1(net253965), .B2(n37745), .C1(net254157), .C2(n37742), 
        .A(n5611), .ZN(n5602) );
  OAI222_X1 U3203 ( .A1(n37967), .A2(n35911), .B1(n38315), .B2(n35399), .C1(
        n38143), .C2(n36423), .ZN(n5611) );
  AOI221_X1 U3204 ( .B1(net254189), .B2(n37739), .C1(net253773), .C2(n37736), 
        .A(n5612), .ZN(n5601) );
  OAI222_X1 U3205 ( .A1(n38162), .A2(n35912), .B1(n37979), .B2(n35400), .C1(
        n38338), .C2(n36424), .ZN(n5612) );
  AOI221_X1 U3206 ( .B1(net254093), .B2(n37733), .C1(net254285), .C2(n37730), 
        .A(n5617), .ZN(n5616) );
  OAI222_X1 U3207 ( .A1(n38075), .A2(n35913), .B1(n38423), .B2(n35401), .C1(
        n38251), .C2(n36425), .ZN(n5617) );
  AOI221_X1 U3208 ( .B1(net254317), .B2(n37727), .C1(net253901), .C2(n37724), 
        .A(n5618), .ZN(n5615) );
  OAI222_X1 U3209 ( .A1(n38270), .A2(n35914), .B1(n38087), .B2(n35402), .C1(
        n38446), .C2(n36426), .ZN(n5618) );
  AOI221_X1 U3210 ( .B1(net254253), .B2(n37721), .C1(net253837), .C2(n37718), 
        .A(n5619), .ZN(n5614) );
  OAI222_X1 U3211 ( .A1(n38216), .A2(n35915), .B1(n38033), .B2(n35403), .C1(
        n38392), .C2(n36427), .ZN(n5619) );
  AOI221_X1 U3212 ( .B1(net253869), .B2(n37715), .C1(net254061), .C2(n37712), 
        .A(n5620), .ZN(n5613) );
  OAI222_X1 U3213 ( .A1(n38411), .A2(n35916), .B1(n38228), .B2(n35404), .C1(
        n38056), .C2(n36428), .ZN(n5620) );
  AOI221_X1 U3214 ( .B1(net253678), .B2(n37784), .C1(net253646), .C2(n37781), 
        .A(n5524), .ZN(n5521) );
  OAI222_X1 U3215 ( .A1(n37838), .A2(n35917), .B1(n37814), .B2(n35405), .C1(
        n37828), .C2(n36429), .ZN(n5524) );
  AOI221_X1 U3216 ( .B1(net253806), .B2(n37757), .C1(net253998), .C2(n37754), 
        .A(n5549), .ZN(n5546) );
  OAI222_X1 U3217 ( .A1(n38357), .A2(n35918), .B1(n38174), .B2(n35406), .C1(
        n38002), .C2(n36430), .ZN(n5549) );
  AOI221_X1 U3218 ( .B1(net254030), .B2(n37751), .C1(net254222), .C2(n37748), 
        .A(n5552), .ZN(n5545) );
  OAI222_X1 U3219 ( .A1(n38021), .A2(n35919), .B1(n38369), .B2(n35407), .C1(
        n38197), .C2(n36431), .ZN(n5552) );
  AOI221_X1 U3220 ( .B1(net253966), .B2(n37745), .C1(net254158), .C2(n37742), 
        .A(n5557), .ZN(n5544) );
  OAI222_X1 U3221 ( .A1(n37967), .A2(n35920), .B1(n38315), .B2(n35408), .C1(
        n38143), .C2(n36432), .ZN(n5557) );
  AOI221_X1 U3222 ( .B1(net254190), .B2(n37739), .C1(net253774), .C2(n37736), 
        .A(n5562), .ZN(n5543) );
  OAI222_X1 U3223 ( .A1(n38162), .A2(n35921), .B1(n37979), .B2(n35409), .C1(
        n38338), .C2(n36433), .ZN(n5562) );
  AOI221_X1 U3224 ( .B1(net254094), .B2(n37733), .C1(net254286), .C2(n37730), 
        .A(n5569), .ZN(n5566) );
  OAI222_X1 U3225 ( .A1(n38075), .A2(n35922), .B1(n38423), .B2(n35410), .C1(
        n38251), .C2(n36434), .ZN(n5569) );
  AOI221_X1 U3226 ( .B1(net254318), .B2(n37727), .C1(net253902), .C2(n37724), 
        .A(n5572), .ZN(n5565) );
  OAI222_X1 U3227 ( .A1(n38270), .A2(n35923), .B1(n38087), .B2(n35411), .C1(
        n38446), .C2(n36435), .ZN(n5572) );
  AOI221_X1 U3228 ( .B1(net254254), .B2(n37721), .C1(net253838), .C2(n37718), 
        .A(n5575), .ZN(n5564) );
  OAI222_X1 U3229 ( .A1(n38216), .A2(n35924), .B1(n38033), .B2(n35412), .C1(
        n38392), .C2(n36436), .ZN(n5575) );
  AOI221_X1 U3230 ( .B1(net253870), .B2(n37715), .C1(net254062), .C2(n37712), 
        .A(n5578), .ZN(n5563) );
  OAI222_X1 U3231 ( .A1(n38411), .A2(n35925), .B1(n38228), .B2(n35413), .C1(
        n38056), .C2(n36437), .ZN(n5578) );
  AOI221_X1 U3232 ( .B1(net253647), .B2(n37782), .C1(net253615), .C2(n37779), 
        .A(n9570), .ZN(n9569) );
  OAI222_X1 U3233 ( .A1(n37840), .A2(n35926), .B1(n37816), .B2(n35414), .C1(
        n37826), .C2(n36438), .ZN(n9570) );
  AOI221_X1 U3234 ( .B1(n38617), .B2(n6368), .C1(n38605), .C2(n9602), .A(n9596), .ZN(n9595) );
  OAI222_X1 U3235 ( .A1(n38593), .A2(n35927), .B1(n38569), .B2(n35415), .C1(
        n38579), .C2(n36439), .ZN(n9596) );
  AOI221_X1 U3236 ( .B1(net253775), .B2(n37755), .C1(net253967), .C2(n37752), 
        .A(n9612), .ZN(n9611) );
  OAI222_X1 U3237 ( .A1(n38359), .A2(n35928), .B1(n38176), .B2(n35416), .C1(
        n38000), .C2(n36440), .ZN(n9612) );
  AOI221_X1 U3238 ( .B1(net254063), .B2(n37731), .C1(net254255), .C2(n37728), 
        .A(n9624), .ZN(n9623) );
  OAI222_X1 U3239 ( .A1(n38077), .A2(n35929), .B1(n38425), .B2(n35417), .C1(
        n38249), .C2(n36441), .ZN(n9624) );
  AOI221_X1 U3240 ( .B1(net253648), .B2(n37782), .C1(net253616), .C2(n37779), 
        .A(n9527), .ZN(n9526) );
  OAI222_X1 U3241 ( .A1(n37840), .A2(n35930), .B1(n37816), .B2(n35418), .C1(
        n37826), .C2(n36442), .ZN(n9527) );
  AOI221_X1 U3242 ( .B1(n38617), .B2(n6369), .C1(n38605), .C2(n9542), .A(n9535), .ZN(n9534) );
  OAI222_X1 U3243 ( .A1(n38593), .A2(n35931), .B1(n38569), .B2(n35419), .C1(
        n38579), .C2(n36443), .ZN(n9535) );
  AOI221_X1 U3244 ( .B1(net253776), .B2(n37755), .C1(net253968), .C2(n37752), 
        .A(n9545), .ZN(n9543) );
  OAI222_X1 U3245 ( .A1(n38359), .A2(n35932), .B1(n38176), .B2(n35420), .C1(
        n38000), .C2(n36444), .ZN(n9545) );
  AOI221_X1 U3246 ( .B1(net254064), .B2(n37731), .C1(net254256), .C2(n37728), 
        .A(n9555), .ZN(n9554) );
  OAI222_X1 U3247 ( .A1(n38077), .A2(n35933), .B1(n38425), .B2(n35421), .C1(
        n38249), .C2(n36445), .ZN(n9555) );
  AOI221_X1 U3248 ( .B1(net253649), .B2(n37782), .C1(net253617), .C2(n37779), 
        .A(n9485), .ZN(n9484) );
  OAI222_X1 U3249 ( .A1(n37840), .A2(n35934), .B1(n37816), .B2(n35422), .C1(
        n37826), .C2(n36446), .ZN(n9485) );
  AOI221_X1 U3250 ( .B1(n38617), .B2(n6370), .C1(n38605), .C2(n9500), .A(n9493), .ZN(n9492) );
  OAI222_X1 U3251 ( .A1(n38593), .A2(n35935), .B1(n38569), .B2(n35423), .C1(
        n38579), .C2(n36447), .ZN(n9493) );
  AOI221_X1 U3252 ( .B1(net253777), .B2(n37755), .C1(net253969), .C2(n37752), 
        .A(n9503), .ZN(n9501) );
  OAI222_X1 U3253 ( .A1(n38359), .A2(n35936), .B1(n38176), .B2(n35424), .C1(
        n38000), .C2(n36448), .ZN(n9503) );
  AOI221_X1 U3254 ( .B1(net254065), .B2(n37731), .C1(net254257), .C2(n37728), 
        .A(n9513), .ZN(n9512) );
  OAI222_X1 U3255 ( .A1(n38077), .A2(n35937), .B1(n38425), .B2(n35425), .C1(
        n38249), .C2(n36449), .ZN(n9513) );
  AOI221_X1 U3256 ( .B1(net253650), .B2(n37782), .C1(net253618), .C2(n37779), 
        .A(n9443), .ZN(n9442) );
  OAI222_X1 U3257 ( .A1(n37840), .A2(n35938), .B1(n37816), .B2(n35426), .C1(
        n37826), .C2(n36450), .ZN(n9443) );
  AOI221_X1 U3258 ( .B1(n38617), .B2(n6372), .C1(n38605), .C2(n9458), .A(n9451), .ZN(n9450) );
  OAI222_X1 U3259 ( .A1(n38593), .A2(n35939), .B1(n38569), .B2(n35427), .C1(
        n38579), .C2(n36451), .ZN(n9451) );
  AOI221_X1 U3260 ( .B1(net253778), .B2(n37755), .C1(net253970), .C2(n37752), 
        .A(n9461), .ZN(n9459) );
  OAI222_X1 U3261 ( .A1(n38359), .A2(n35940), .B1(n38176), .B2(n35428), .C1(
        n38000), .C2(n36452), .ZN(n9461) );
  AOI221_X1 U3262 ( .B1(net254066), .B2(n37731), .C1(net254258), .C2(n37728), 
        .A(n9471), .ZN(n9470) );
  OAI222_X1 U3263 ( .A1(n38077), .A2(n35941), .B1(n38425), .B2(n35429), .C1(
        n38249), .C2(n36453), .ZN(n9471) );
  AOI221_X1 U3264 ( .B1(net253651), .B2(n37782), .C1(net253619), .C2(n37779), 
        .A(n9401), .ZN(n9400) );
  OAI222_X1 U3265 ( .A1(n37840), .A2(n35942), .B1(n37816), .B2(n35430), .C1(
        n37826), .C2(n36454), .ZN(n9401) );
  AOI221_X1 U3266 ( .B1(n38617), .B2(n6374), .C1(n38605), .C2(n9416), .A(n9409), .ZN(n9408) );
  OAI222_X1 U3267 ( .A1(n38593), .A2(n35943), .B1(n38569), .B2(n35431), .C1(
        n38579), .C2(n36455), .ZN(n9409) );
  AOI221_X1 U3268 ( .B1(net253779), .B2(n37755), .C1(net253971), .C2(n37752), 
        .A(n9419), .ZN(n9417) );
  OAI222_X1 U3269 ( .A1(n38359), .A2(n35944), .B1(n38176), .B2(n35432), .C1(
        n38000), .C2(n36456), .ZN(n9419) );
  AOI221_X1 U3270 ( .B1(net254067), .B2(n37731), .C1(net254259), .C2(n37728), 
        .A(n9429), .ZN(n9428) );
  OAI222_X1 U3271 ( .A1(n38077), .A2(n35945), .B1(n38425), .B2(n35433), .C1(
        n38249), .C2(n36457), .ZN(n9429) );
  AOI221_X1 U3272 ( .B1(net253652), .B2(n37782), .C1(net253620), .C2(n37779), 
        .A(n9359), .ZN(n9358) );
  OAI222_X1 U3273 ( .A1(n37840), .A2(n35946), .B1(n37816), .B2(n35434), .C1(
        n37826), .C2(n36458), .ZN(n9359) );
  AOI221_X1 U3274 ( .B1(n38617), .B2(n6375), .C1(n38605), .C2(n9374), .A(n9367), .ZN(n9366) );
  OAI222_X1 U3275 ( .A1(n38593), .A2(n35947), .B1(n38569), .B2(n35435), .C1(
        n38579), .C2(n36459), .ZN(n9367) );
  AOI221_X1 U3276 ( .B1(net253780), .B2(n37755), .C1(net253972), .C2(n37752), 
        .A(n9377), .ZN(n9375) );
  OAI222_X1 U3277 ( .A1(n38359), .A2(n35948), .B1(n38176), .B2(n35436), .C1(
        n38000), .C2(n36460), .ZN(n9377) );
  AOI221_X1 U3278 ( .B1(net254068), .B2(n37731), .C1(net254260), .C2(n37728), 
        .A(n9387), .ZN(n9386) );
  OAI222_X1 U3279 ( .A1(n38077), .A2(n35949), .B1(n38425), .B2(n35437), .C1(
        n38249), .C2(n36461), .ZN(n9387) );
  AOI221_X1 U3280 ( .B1(net253653), .B2(n37782), .C1(net253621), .C2(n37779), 
        .A(n9317), .ZN(n9316) );
  OAI222_X1 U3281 ( .A1(n37840), .A2(n35950), .B1(n37816), .B2(n35438), .C1(
        n37826), .C2(n36462), .ZN(n9317) );
  AOI221_X1 U3282 ( .B1(n38617), .B2(n6376), .C1(n38605), .C2(n9332), .A(n9325), .ZN(n9324) );
  OAI222_X1 U3283 ( .A1(n38593), .A2(n35951), .B1(n38569), .B2(n35439), .C1(
        n38579), .C2(n36463), .ZN(n9325) );
  AOI221_X1 U3284 ( .B1(net253781), .B2(n37755), .C1(net253973), .C2(n37752), 
        .A(n9335), .ZN(n9333) );
  OAI222_X1 U3285 ( .A1(n38359), .A2(n35952), .B1(n38176), .B2(n35440), .C1(
        n38000), .C2(n36464), .ZN(n9335) );
  AOI221_X1 U3286 ( .B1(net254069), .B2(n37731), .C1(net254261), .C2(n37728), 
        .A(n9345), .ZN(n9344) );
  OAI222_X1 U3287 ( .A1(n38077), .A2(n35953), .B1(n38425), .B2(n35441), .C1(
        n38249), .C2(n36465), .ZN(n9345) );
  AOI221_X1 U3288 ( .B1(net253654), .B2(n37782), .C1(net253622), .C2(n37779), 
        .A(n9275), .ZN(n9274) );
  OAI222_X1 U3289 ( .A1(n37840), .A2(n35954), .B1(n37816), .B2(n35442), .C1(
        n37826), .C2(n36466), .ZN(n9275) );
  AOI221_X1 U3290 ( .B1(n38617), .B2(n6377), .C1(n38604), .C2(n9290), .A(n9283), .ZN(n9282) );
  OAI222_X1 U3291 ( .A1(n38593), .A2(n35955), .B1(n38569), .B2(n35443), .C1(
        n38579), .C2(n36467), .ZN(n9283) );
  AOI221_X1 U3292 ( .B1(net253782), .B2(n37755), .C1(net253974), .C2(n37752), 
        .A(n9293), .ZN(n9291) );
  OAI222_X1 U3293 ( .A1(n38359), .A2(n35956), .B1(n38176), .B2(n35444), .C1(
        n38000), .C2(n36468), .ZN(n9293) );
  AOI221_X1 U3294 ( .B1(net254070), .B2(n37731), .C1(net254262), .C2(n37728), 
        .A(n9303), .ZN(n9302) );
  OAI222_X1 U3295 ( .A1(n38077), .A2(n35957), .B1(n38425), .B2(n35445), .C1(
        n38249), .C2(n36469), .ZN(n9303) );
  AOI221_X1 U3296 ( .B1(net253655), .B2(n37782), .C1(net253623), .C2(n37779), 
        .A(n6641), .ZN(n6640) );
  OAI222_X1 U3297 ( .A1(n37840), .A2(n35958), .B1(n37816), .B2(n35446), .C1(
        n37826), .C2(n36470), .ZN(n6641) );
  AOI221_X1 U3298 ( .B1(n38617), .B2(n6378), .C1(n38604), .C2(n6656), .A(n6649), .ZN(n6648) );
  OAI222_X1 U3299 ( .A1(n38593), .A2(n35959), .B1(n38569), .B2(n35447), .C1(
        n38579), .C2(n36471), .ZN(n6649) );
  AOI221_X1 U3300 ( .B1(net253783), .B2(n37755), .C1(net253975), .C2(n37752), 
        .A(n6659), .ZN(n6657) );
  OAI222_X1 U3301 ( .A1(n38359), .A2(n35960), .B1(n38176), .B2(n35448), .C1(
        n38000), .C2(n36472), .ZN(n6659) );
  AOI221_X1 U3302 ( .B1(net254071), .B2(n37731), .C1(net254263), .C2(n37728), 
        .A(n6669), .ZN(n6668) );
  OAI222_X1 U3303 ( .A1(n38077), .A2(n35961), .B1(n38425), .B2(n35449), .C1(
        n38249), .C2(n36473), .ZN(n6669) );
  AOI221_X1 U3304 ( .B1(net253656), .B2(n37782), .C1(net253624), .C2(n37779), 
        .A(n6599), .ZN(n6598) );
  OAI222_X1 U3305 ( .A1(n37839), .A2(n35962), .B1(n37815), .B2(n35450), .C1(
        n37826), .C2(n36474), .ZN(n6599) );
  AOI221_X1 U3306 ( .B1(n38616), .B2(n6379), .C1(n38604), .C2(n6614), .A(n6607), .ZN(n6606) );
  OAI222_X1 U3307 ( .A1(n38592), .A2(n35963), .B1(n38568), .B2(n35451), .C1(
        n38579), .C2(n36475), .ZN(n6607) );
  AOI221_X1 U3308 ( .B1(net253784), .B2(n37755), .C1(net253976), .C2(n37752), 
        .A(n6617), .ZN(n6615) );
  OAI222_X1 U3309 ( .A1(n38358), .A2(n35964), .B1(n38175), .B2(n35452), .C1(
        n38000), .C2(n36476), .ZN(n6617) );
  AOI221_X1 U3310 ( .B1(net254072), .B2(n37731), .C1(net254264), .C2(n37728), 
        .A(n6627), .ZN(n6626) );
  OAI222_X1 U3311 ( .A1(n38076), .A2(n35965), .B1(n38424), .B2(n35453), .C1(
        n38249), .C2(n36477), .ZN(n6627) );
  AOI221_X1 U3312 ( .B1(net253657), .B2(n37782), .C1(net253625), .C2(n37779), 
        .A(n6557), .ZN(n6556) );
  OAI222_X1 U3313 ( .A1(n37839), .A2(n35966), .B1(n37815), .B2(n35454), .C1(
        n37826), .C2(n36478), .ZN(n6557) );
  AOI221_X1 U3314 ( .B1(n38616), .B2(n6380), .C1(n38604), .C2(n6572), .A(n6565), .ZN(n6564) );
  OAI222_X1 U3315 ( .A1(n38592), .A2(n35967), .B1(n38568), .B2(n35455), .C1(
        n38579), .C2(n36479), .ZN(n6565) );
  AOI221_X1 U3316 ( .B1(net253785), .B2(n37755), .C1(net253977), .C2(n37752), 
        .A(n6575), .ZN(n6573) );
  OAI222_X1 U3317 ( .A1(n38358), .A2(n35968), .B1(n38175), .B2(n35456), .C1(
        n38000), .C2(n36480), .ZN(n6575) );
  AOI221_X1 U3318 ( .B1(net254073), .B2(n37731), .C1(net254265), .C2(n37728), 
        .A(n6585), .ZN(n6584) );
  OAI222_X1 U3319 ( .A1(n38076), .A2(n35969), .B1(n38424), .B2(n35457), .C1(
        n38249), .C2(n36481), .ZN(n6585) );
  AOI221_X1 U3320 ( .B1(net253658), .B2(n37782), .C1(net253626), .C2(n37779), 
        .A(n6515), .ZN(n6514) );
  OAI222_X1 U3321 ( .A1(n37839), .A2(n35970), .B1(n37815), .B2(n35458), .C1(
        n37826), .C2(n36482), .ZN(n6515) );
  AOI221_X1 U3322 ( .B1(n38616), .B2(n6381), .C1(n38604), .C2(n6530), .A(n6523), .ZN(n6522) );
  OAI222_X1 U3323 ( .A1(n38592), .A2(n35971), .B1(n38568), .B2(n35459), .C1(
        n38579), .C2(n36483), .ZN(n6523) );
  AOI221_X1 U3324 ( .B1(net253786), .B2(n37755), .C1(net253978), .C2(n37752), 
        .A(n6533), .ZN(n6531) );
  OAI222_X1 U3325 ( .A1(n38358), .A2(n35972), .B1(n38175), .B2(n35460), .C1(
        n38000), .C2(n36484), .ZN(n6533) );
  AOI221_X1 U3326 ( .B1(net254074), .B2(n37731), .C1(net254266), .C2(n37728), 
        .A(n6543), .ZN(n6542) );
  OAI222_X1 U3327 ( .A1(n38076), .A2(n35973), .B1(n38424), .B2(n35461), .C1(
        n38249), .C2(n36485), .ZN(n6543) );
  AOI221_X1 U3328 ( .B1(net253659), .B2(n37783), .C1(net253627), .C2(n37780), 
        .A(n6345), .ZN(n6344) );
  OAI222_X1 U3329 ( .A1(n37839), .A2(n35974), .B1(n37815), .B2(n35462), .C1(
        n37827), .C2(n36486), .ZN(n6345) );
  AOI221_X1 U3330 ( .B1(n38616), .B2(n6382), .C1(n38604), .C2(n6360), .A(n6353), .ZN(n6352) );
  OAI222_X1 U3331 ( .A1(n38592), .A2(n35975), .B1(n38568), .B2(n35463), .C1(
        n38580), .C2(n36487), .ZN(n6353) );
  AOI221_X1 U3332 ( .B1(net253787), .B2(n37756), .C1(net253979), .C2(n37753), 
        .A(n6363), .ZN(n6361) );
  OAI222_X1 U3333 ( .A1(n38358), .A2(n35976), .B1(n38175), .B2(n35464), .C1(
        n38001), .C2(n36488), .ZN(n6363) );
  AOI221_X1 U3334 ( .B1(net254075), .B2(n37732), .C1(net254267), .C2(n37729), 
        .A(n6443), .ZN(n6441) );
  OAI222_X1 U3335 ( .A1(n38076), .A2(n35977), .B1(n38424), .B2(n35465), .C1(
        n38250), .C2(n36489), .ZN(n6443) );
  AOI221_X1 U3336 ( .B1(net253660), .B2(n37783), .C1(net253628), .C2(n37780), 
        .A(n6303), .ZN(n6302) );
  OAI222_X1 U3337 ( .A1(n37839), .A2(n35978), .B1(n37815), .B2(n35466), .C1(
        n37827), .C2(n36490), .ZN(n6303) );
  AOI221_X1 U3338 ( .B1(n38616), .B2(n6383), .C1(n38604), .C2(n6318), .A(n6311), .ZN(n6310) );
  OAI222_X1 U3339 ( .A1(n38592), .A2(n35979), .B1(n38568), .B2(n35467), .C1(
        n38580), .C2(n36491), .ZN(n6311) );
  AOI221_X1 U3340 ( .B1(net253788), .B2(n37756), .C1(net253980), .C2(n37753), 
        .A(n6321), .ZN(n6319) );
  OAI222_X1 U3341 ( .A1(n38358), .A2(n35980), .B1(n38175), .B2(n35468), .C1(
        n38001), .C2(n36492), .ZN(n6321) );
  AOI221_X1 U3342 ( .B1(net254076), .B2(n37732), .C1(net254268), .C2(n37729), 
        .A(n6331), .ZN(n6330) );
  OAI222_X1 U3343 ( .A1(n38076), .A2(n35981), .B1(n38424), .B2(n35469), .C1(
        n38250), .C2(n36493), .ZN(n6331) );
  AOI221_X1 U3344 ( .B1(net253661), .B2(n37783), .C1(net253629), .C2(n37780), 
        .A(n6261), .ZN(n6260) );
  OAI222_X1 U3345 ( .A1(n37839), .A2(n35982), .B1(n37815), .B2(n35470), .C1(
        n37827), .C2(n36494), .ZN(n6261) );
  AOI221_X1 U3346 ( .B1(n38616), .B2(n6384), .C1(n38604), .C2(n6276), .A(n6269), .ZN(n6268) );
  OAI222_X1 U3347 ( .A1(n38592), .A2(n35983), .B1(n38568), .B2(n35471), .C1(
        n38580), .C2(n36495), .ZN(n6269) );
  AOI221_X1 U3348 ( .B1(net253789), .B2(n37756), .C1(net253981), .C2(n37753), 
        .A(n6279), .ZN(n6277) );
  OAI222_X1 U3349 ( .A1(n38358), .A2(n35984), .B1(n38175), .B2(n35472), .C1(
        n38001), .C2(n36496), .ZN(n6279) );
  AOI221_X1 U3350 ( .B1(net254077), .B2(n37732), .C1(net254269), .C2(n37729), 
        .A(n6289), .ZN(n6288) );
  OAI222_X1 U3351 ( .A1(n38076), .A2(n35985), .B1(n38424), .B2(n35473), .C1(
        n38250), .C2(n36497), .ZN(n6289) );
  AOI221_X1 U3352 ( .B1(net253662), .B2(n37783), .C1(net253630), .C2(n37780), 
        .A(n6219), .ZN(n6218) );
  OAI222_X1 U3353 ( .A1(n37839), .A2(n35986), .B1(n37815), .B2(n35474), .C1(
        n37827), .C2(n36498), .ZN(n6219) );
  AOI221_X1 U3354 ( .B1(n38616), .B2(n6385), .C1(n38604), .C2(n6234), .A(n6227), .ZN(n6226) );
  OAI222_X1 U3355 ( .A1(n38592), .A2(n35987), .B1(n38568), .B2(n35475), .C1(
        n38580), .C2(n36499), .ZN(n6227) );
  AOI221_X1 U3356 ( .B1(net253790), .B2(n37756), .C1(net253982), .C2(n37753), 
        .A(n6237), .ZN(n6235) );
  OAI222_X1 U3357 ( .A1(n38358), .A2(n35988), .B1(n38175), .B2(n35476), .C1(
        n38001), .C2(n36500), .ZN(n6237) );
  AOI221_X1 U3358 ( .B1(net254078), .B2(n37732), .C1(net254270), .C2(n37729), 
        .A(n6247), .ZN(n6246) );
  OAI222_X1 U3359 ( .A1(n38076), .A2(n35989), .B1(n38424), .B2(n35477), .C1(
        n38250), .C2(n36501), .ZN(n6247) );
  AOI221_X1 U3360 ( .B1(net253663), .B2(n37783), .C1(net253631), .C2(n37780), 
        .A(n6177), .ZN(n6176) );
  OAI222_X1 U3361 ( .A1(n37839), .A2(n35990), .B1(n37815), .B2(n35478), .C1(
        n37827), .C2(n36502), .ZN(n6177) );
  AOI221_X1 U3362 ( .B1(n38616), .B2(n6386), .C1(n38604), .C2(n6192), .A(n6185), .ZN(n6184) );
  OAI222_X1 U3363 ( .A1(n38592), .A2(n35991), .B1(n38568), .B2(n35479), .C1(
        n38580), .C2(n36503), .ZN(n6185) );
  AOI221_X1 U3364 ( .B1(net253791), .B2(n37756), .C1(net253983), .C2(n37753), 
        .A(n6195), .ZN(n6193) );
  OAI222_X1 U3365 ( .A1(n38358), .A2(n35992), .B1(n38175), .B2(n35480), .C1(
        n38001), .C2(n36504), .ZN(n6195) );
  AOI221_X1 U3366 ( .B1(net254079), .B2(n37732), .C1(net254271), .C2(n37729), 
        .A(n6205), .ZN(n6204) );
  OAI222_X1 U3367 ( .A1(n38076), .A2(n35993), .B1(n38424), .B2(n35481), .C1(
        n38250), .C2(n36505), .ZN(n6205) );
  AOI221_X1 U3368 ( .B1(net253664), .B2(n37783), .C1(net253632), .C2(n37780), 
        .A(n6135), .ZN(n6134) );
  OAI222_X1 U3369 ( .A1(n37839), .A2(n35994), .B1(n37815), .B2(n35482), .C1(
        n37827), .C2(n36506), .ZN(n6135) );
  AOI221_X1 U3370 ( .B1(n38616), .B2(n6387), .C1(n38604), .C2(n6150), .A(n6143), .ZN(n6142) );
  OAI222_X1 U3371 ( .A1(n38592), .A2(n35995), .B1(n38568), .B2(n35483), .C1(
        n38580), .C2(n36507), .ZN(n6143) );
  AOI221_X1 U3372 ( .B1(net253792), .B2(n37756), .C1(net253984), .C2(n37753), 
        .A(n6153), .ZN(n6151) );
  OAI222_X1 U3373 ( .A1(n38358), .A2(n35996), .B1(n38175), .B2(n35484), .C1(
        n38001), .C2(n36508), .ZN(n6153) );
  AOI221_X1 U3374 ( .B1(net254080), .B2(n37732), .C1(net254272), .C2(n37729), 
        .A(n6163), .ZN(n6162) );
  OAI222_X1 U3375 ( .A1(n38076), .A2(n35997), .B1(n38424), .B2(n35485), .C1(
        n38250), .C2(n36509), .ZN(n6163) );
  AOI221_X1 U3376 ( .B1(net253665), .B2(n37783), .C1(net253633), .C2(n37780), 
        .A(n6093), .ZN(n6092) );
  OAI222_X1 U3377 ( .A1(n37839), .A2(n35998), .B1(n37815), .B2(n35486), .C1(
        n37827), .C2(n36510), .ZN(n6093) );
  AOI221_X1 U3378 ( .B1(n38616), .B2(n6388), .C1(n38604), .C2(n6108), .A(n6101), .ZN(n6100) );
  OAI222_X1 U3379 ( .A1(n38592), .A2(n35999), .B1(n38568), .B2(n35487), .C1(
        n38580), .C2(n36511), .ZN(n6101) );
  AOI221_X1 U3380 ( .B1(net253793), .B2(n37756), .C1(net253985), .C2(n37753), 
        .A(n6111), .ZN(n6109) );
  OAI222_X1 U3381 ( .A1(n38358), .A2(n36000), .B1(n38175), .B2(n35488), .C1(
        n38001), .C2(n36512), .ZN(n6111) );
  AOI221_X1 U3382 ( .B1(net254081), .B2(n37732), .C1(net254273), .C2(n37729), 
        .A(n6121), .ZN(n6120) );
  OAI222_X1 U3383 ( .A1(n38076), .A2(n36001), .B1(n38424), .B2(n35489), .C1(
        n38250), .C2(n36513), .ZN(n6121) );
  AOI221_X1 U3384 ( .B1(net253666), .B2(n37783), .C1(net253634), .C2(n37780), 
        .A(n6051), .ZN(n6050) );
  OAI222_X1 U3385 ( .A1(n37839), .A2(n36002), .B1(n37815), .B2(n35490), .C1(
        n37827), .C2(n36514), .ZN(n6051) );
  AOI221_X1 U3386 ( .B1(n38616), .B2(n6389), .C1(n38604), .C2(n6066), .A(n6059), .ZN(n6058) );
  OAI222_X1 U3387 ( .A1(n38592), .A2(n36003), .B1(n38568), .B2(n35491), .C1(
        n38580), .C2(n36515), .ZN(n6059) );
  AOI221_X1 U3388 ( .B1(net253794), .B2(n37756), .C1(net253986), .C2(n37753), 
        .A(n6069), .ZN(n6067) );
  OAI222_X1 U3389 ( .A1(n38358), .A2(n36004), .B1(n38175), .B2(n35492), .C1(
        n38001), .C2(n36516), .ZN(n6069) );
  AOI221_X1 U3390 ( .B1(net254082), .B2(n37732), .C1(net254274), .C2(n37729), 
        .A(n6079), .ZN(n6078) );
  OAI222_X1 U3391 ( .A1(n38076), .A2(n36005), .B1(n38424), .B2(n35493), .C1(
        n38250), .C2(n36517), .ZN(n6079) );
  AOI221_X1 U3392 ( .B1(net253667), .B2(n37783), .C1(net253635), .C2(n37780), 
        .A(n6009), .ZN(n6008) );
  OAI222_X1 U3393 ( .A1(n37839), .A2(n36006), .B1(n37815), .B2(n35494), .C1(
        n37827), .C2(n36518), .ZN(n6009) );
  AOI221_X1 U3394 ( .B1(n38616), .B2(n6390), .C1(n38603), .C2(n6024), .A(n6017), .ZN(n6016) );
  OAI222_X1 U3395 ( .A1(n38592), .A2(n36007), .B1(n38568), .B2(n35495), .C1(
        n38580), .C2(n36519), .ZN(n6017) );
  AOI221_X1 U3396 ( .B1(net253795), .B2(n37756), .C1(net253987), .C2(n37753), 
        .A(n6027), .ZN(n6025) );
  OAI222_X1 U3397 ( .A1(n38358), .A2(n36008), .B1(n38175), .B2(n35496), .C1(
        n38001), .C2(n36520), .ZN(n6027) );
  AOI221_X1 U3398 ( .B1(net254083), .B2(n37732), .C1(net254275), .C2(n37729), 
        .A(n6037), .ZN(n6036) );
  OAI222_X1 U3399 ( .A1(n38076), .A2(n36009), .B1(n38424), .B2(n35497), .C1(
        n38250), .C2(n36521), .ZN(n6037) );
  AOI221_X1 U3400 ( .B1(net253668), .B2(n37783), .C1(net253636), .C2(n37780), 
        .A(n5967), .ZN(n5966) );
  OAI222_X1 U3401 ( .A1(n37838), .A2(n36010), .B1(n37814), .B2(n35498), .C1(
        n37827), .C2(n36522), .ZN(n5967) );
  AOI221_X1 U3402 ( .B1(n38615), .B2(n6391), .C1(n38603), .C2(n5982), .A(n5975), .ZN(n5974) );
  OAI222_X1 U3403 ( .A1(n38591), .A2(n36011), .B1(n38567), .B2(n35499), .C1(
        n38580), .C2(n36523), .ZN(n5975) );
  AOI221_X1 U3404 ( .B1(net253796), .B2(n37756), .C1(net253988), .C2(n37753), 
        .A(n5985), .ZN(n5983) );
  OAI222_X1 U3405 ( .A1(n38357), .A2(n36012), .B1(n38174), .B2(n35500), .C1(
        n38001), .C2(n36524), .ZN(n5985) );
  AOI221_X1 U3406 ( .B1(net254084), .B2(n37732), .C1(net254276), .C2(n37729), 
        .A(n5995), .ZN(n5994) );
  OAI222_X1 U3407 ( .A1(n38075), .A2(n36013), .B1(n38423), .B2(n35501), .C1(
        n38250), .C2(n36525), .ZN(n5995) );
  AOI221_X1 U3408 ( .B1(net253669), .B2(n37783), .C1(net253637), .C2(n37780), 
        .A(n5925), .ZN(n5924) );
  OAI222_X1 U3409 ( .A1(n37838), .A2(n36014), .B1(n37814), .B2(n35502), .C1(
        n37827), .C2(n36526), .ZN(n5925) );
  AOI221_X1 U3410 ( .B1(n38615), .B2(n6392), .C1(n38603), .C2(n5940), .A(n5933), .ZN(n5932) );
  OAI222_X1 U3411 ( .A1(n38591), .A2(n36015), .B1(n38567), .B2(n35503), .C1(
        n38580), .C2(n36527), .ZN(n5933) );
  AOI221_X1 U3412 ( .B1(net253797), .B2(n37756), .C1(net253989), .C2(n37753), 
        .A(n5943), .ZN(n5941) );
  OAI222_X1 U3413 ( .A1(n38357), .A2(n36016), .B1(n38174), .B2(n35504), .C1(
        n38001), .C2(n36528), .ZN(n5943) );
  AOI221_X1 U3414 ( .B1(net254085), .B2(n37732), .C1(net254277), .C2(n37729), 
        .A(n5953), .ZN(n5952) );
  OAI222_X1 U3415 ( .A1(n38075), .A2(n36017), .B1(n38423), .B2(n35505), .C1(
        n38250), .C2(n36529), .ZN(n5953) );
  AOI221_X1 U3416 ( .B1(net253670), .B2(n37783), .C1(net253638), .C2(n37780), 
        .A(n5883), .ZN(n5882) );
  OAI222_X1 U3417 ( .A1(n37838), .A2(n36018), .B1(n37814), .B2(n35506), .C1(
        n37827), .C2(n36530), .ZN(n5883) );
  AOI221_X1 U3418 ( .B1(n38615), .B2(n6393), .C1(n38603), .C2(n5898), .A(n5891), .ZN(n5890) );
  OAI222_X1 U3419 ( .A1(n38591), .A2(n36019), .B1(n38567), .B2(n35507), .C1(
        n38580), .C2(n36531), .ZN(n5891) );
  AOI221_X1 U3420 ( .B1(net253798), .B2(n37756), .C1(net253990), .C2(n37753), 
        .A(n5901), .ZN(n5899) );
  OAI222_X1 U3421 ( .A1(n38357), .A2(n36020), .B1(n38174), .B2(n35508), .C1(
        n38001), .C2(n36532), .ZN(n5901) );
  AOI221_X1 U3422 ( .B1(net254086), .B2(n37732), .C1(net254278), .C2(n37729), 
        .A(n5911), .ZN(n5910) );
  OAI222_X1 U3423 ( .A1(n38075), .A2(n36021), .B1(n38423), .B2(n35509), .C1(
        n38250), .C2(n36533), .ZN(n5911) );
  AOI221_X1 U3424 ( .B1(n38615), .B2(n6394), .C1(n38603), .C2(n5856), .A(n5849), .ZN(n5848) );
  OAI222_X1 U3425 ( .A1(n38591), .A2(n36022), .B1(n38567), .B2(n35510), .C1(
        n38581), .C2(n36534), .ZN(n5849) );
  AOI221_X1 U3426 ( .B1(n38615), .B2(n6395), .C1(n38603), .C2(n5814), .A(n5807), .ZN(n5806) );
  OAI222_X1 U3427 ( .A1(n38591), .A2(n36023), .B1(n38567), .B2(n35511), .C1(
        n38581), .C2(n36535), .ZN(n5807) );
  AOI221_X1 U3428 ( .B1(n38615), .B2(n6396), .C1(n38603), .C2(n5772), .A(n5765), .ZN(n5764) );
  OAI222_X1 U3429 ( .A1(n38591), .A2(n36024), .B1(n38567), .B2(n35512), .C1(
        n38581), .C2(n36536), .ZN(n5765) );
  AOI221_X1 U3430 ( .B1(n38615), .B2(n6397), .C1(n38603), .C2(n5730), .A(n5723), .ZN(n5722) );
  OAI222_X1 U3431 ( .A1(n38591), .A2(n36025), .B1(n38567), .B2(n35513), .C1(
        n38581), .C2(n36537), .ZN(n5723) );
  AOI221_X1 U3432 ( .B1(n38615), .B2(n6398), .C1(n38603), .C2(n5688), .A(n5681), .ZN(n5680) );
  OAI222_X1 U3433 ( .A1(n38591), .A2(n36026), .B1(n38567), .B2(n35514), .C1(
        n38581), .C2(n36538), .ZN(n5681) );
  AOI221_X1 U3434 ( .B1(n38615), .B2(n6399), .C1(n38603), .C2(n5646), .A(n5639), .ZN(n5638) );
  OAI222_X1 U3435 ( .A1(n38591), .A2(n36027), .B1(n38567), .B2(n35515), .C1(
        n38581), .C2(n36539), .ZN(n5639) );
  AOI221_X1 U3436 ( .B1(n38615), .B2(n6400), .C1(n38603), .C2(n5604), .A(n5597), .ZN(n5596) );
  OAI222_X1 U3437 ( .A1(n38591), .A2(n36028), .B1(n38567), .B2(n35516), .C1(
        n38581), .C2(n36540), .ZN(n5597) );
  AOI221_X1 U3438 ( .B1(n38615), .B2(n6401), .C1(n38603), .C2(n5553), .A(n5538), .ZN(n5537) );
  OAI222_X1 U3439 ( .A1(n38591), .A2(n36029), .B1(n38567), .B2(n35517), .C1(
        n38581), .C2(n36541), .ZN(n5538) );
  AOI221_X1 U3440 ( .B1(net253999), .B2(n37749), .C1(net254191), .C2(n37746), 
        .A(n9616), .ZN(n9610) );
  OAI222_X1 U3441 ( .A1(n38023), .A2(n36030), .B1(n38371), .B2(n35518), .C1(
        n38195), .C2(n36542), .ZN(n9616) );
  AOI221_X1 U3442 ( .B1(net254287), .B2(n37725), .C1(net253871), .C2(n37722), 
        .A(n9626), .ZN(n9622) );
  OAI222_X1 U3443 ( .A1(n38272), .A2(n36031), .B1(n38089), .B2(n35519), .C1(
        n38444), .C2(n36543), .ZN(n9626) );
  AOI221_X1 U3444 ( .B1(net254000), .B2(n37749), .C1(net254192), .C2(n37746), 
        .A(n9547), .ZN(n9541) );
  OAI222_X1 U3445 ( .A1(n38023), .A2(n36032), .B1(n38371), .B2(n35520), .C1(
        n38195), .C2(n36544), .ZN(n9547) );
  AOI221_X1 U3446 ( .B1(net254288), .B2(n37725), .C1(net253872), .C2(n37722), 
        .A(n9556), .ZN(n9553) );
  OAI222_X1 U3447 ( .A1(n38272), .A2(n36033), .B1(n38089), .B2(n35521), .C1(
        n38444), .C2(n36545), .ZN(n9556) );
  AOI221_X1 U3448 ( .B1(net254001), .B2(n37749), .C1(net254193), .C2(n37746), 
        .A(n9505), .ZN(n9499) );
  OAI222_X1 U3449 ( .A1(n38023), .A2(n36034), .B1(n38371), .B2(n35522), .C1(
        n38195), .C2(n36546), .ZN(n9505) );
  AOI221_X1 U3450 ( .B1(net254289), .B2(n37725), .C1(net253873), .C2(n37722), 
        .A(n9514), .ZN(n9511) );
  OAI222_X1 U3451 ( .A1(n38272), .A2(n36035), .B1(n38089), .B2(n35523), .C1(
        n38444), .C2(n36547), .ZN(n9514) );
  AOI221_X1 U3452 ( .B1(net254002), .B2(n37749), .C1(net254194), .C2(n37746), 
        .A(n9463), .ZN(n9457) );
  OAI222_X1 U3453 ( .A1(n38023), .A2(n36036), .B1(n38371), .B2(n35524), .C1(
        n38195), .C2(n36548), .ZN(n9463) );
  AOI221_X1 U3454 ( .B1(net254290), .B2(n37725), .C1(net253874), .C2(n37722), 
        .A(n9472), .ZN(n9469) );
  OAI222_X1 U3455 ( .A1(n38272), .A2(n36037), .B1(n38089), .B2(n35525), .C1(
        n38444), .C2(n36549), .ZN(n9472) );
  AOI221_X1 U3456 ( .B1(net254003), .B2(n37749), .C1(net254195), .C2(n37746), 
        .A(n9421), .ZN(n9415) );
  OAI222_X1 U3457 ( .A1(n38023), .A2(n36038), .B1(n38371), .B2(n35526), .C1(
        n38195), .C2(n36550), .ZN(n9421) );
  AOI221_X1 U3458 ( .B1(net254291), .B2(n37725), .C1(net253875), .C2(n37722), 
        .A(n9430), .ZN(n9427) );
  OAI222_X1 U3459 ( .A1(n38272), .A2(n36039), .B1(n38089), .B2(n35527), .C1(
        n38444), .C2(n36551), .ZN(n9430) );
  AOI221_X1 U3460 ( .B1(net254004), .B2(n37749), .C1(net254196), .C2(n37746), 
        .A(n9379), .ZN(n9373) );
  OAI222_X1 U3461 ( .A1(n38023), .A2(n36040), .B1(n38371), .B2(n35528), .C1(
        n38195), .C2(n36552), .ZN(n9379) );
  AOI221_X1 U3462 ( .B1(net254292), .B2(n37725), .C1(net253876), .C2(n37722), 
        .A(n9388), .ZN(n9385) );
  OAI222_X1 U3463 ( .A1(n38272), .A2(n36041), .B1(n38089), .B2(n35529), .C1(
        n38444), .C2(n36553), .ZN(n9388) );
  AOI221_X1 U3464 ( .B1(net254005), .B2(n37749), .C1(net254197), .C2(n37746), 
        .A(n9337), .ZN(n9331) );
  OAI222_X1 U3465 ( .A1(n38023), .A2(n36042), .B1(n38371), .B2(n35530), .C1(
        n38195), .C2(n36554), .ZN(n9337) );
  AOI221_X1 U3466 ( .B1(net254293), .B2(n37725), .C1(net253877), .C2(n37722), 
        .A(n9346), .ZN(n9343) );
  OAI222_X1 U3467 ( .A1(n38272), .A2(n36043), .B1(n38089), .B2(n35531), .C1(
        n38444), .C2(n36555), .ZN(n9346) );
  AOI221_X1 U3468 ( .B1(net254006), .B2(n37749), .C1(net254198), .C2(n37746), 
        .A(n9295), .ZN(n9289) );
  OAI222_X1 U3469 ( .A1(n38023), .A2(n36044), .B1(n38371), .B2(n35532), .C1(
        n38195), .C2(n36556), .ZN(n9295) );
  AOI221_X1 U3470 ( .B1(net254294), .B2(n37725), .C1(net253878), .C2(n37722), 
        .A(n9304), .ZN(n9301) );
  OAI222_X1 U3471 ( .A1(n38272), .A2(n36045), .B1(n38089), .B2(n35533), .C1(
        n38444), .C2(n36557), .ZN(n9304) );
  AOI221_X1 U3472 ( .B1(net254007), .B2(n37749), .C1(net254199), .C2(n37746), 
        .A(n6661), .ZN(n6655) );
  OAI222_X1 U3473 ( .A1(n38023), .A2(n36046), .B1(n38371), .B2(n35534), .C1(
        n38195), .C2(n36558), .ZN(n6661) );
  AOI221_X1 U3474 ( .B1(net254295), .B2(n37725), .C1(net253879), .C2(n37722), 
        .A(n6670), .ZN(n6667) );
  OAI222_X1 U3475 ( .A1(n38272), .A2(n36047), .B1(n38089), .B2(n35535), .C1(
        n38444), .C2(n36559), .ZN(n6670) );
  AOI221_X1 U3476 ( .B1(net254008), .B2(n37749), .C1(net254200), .C2(n37746), 
        .A(n6619), .ZN(n6613) );
  OAI222_X1 U3477 ( .A1(n38022), .A2(n36048), .B1(n38370), .B2(n35536), .C1(
        n38195), .C2(n36560), .ZN(n6619) );
  AOI221_X1 U3478 ( .B1(net254296), .B2(n37725), .C1(net253880), .C2(n37722), 
        .A(n6628), .ZN(n6625) );
  OAI222_X1 U3479 ( .A1(n38271), .A2(n36049), .B1(n38088), .B2(n35537), .C1(
        n38444), .C2(n36561), .ZN(n6628) );
  AOI221_X1 U3480 ( .B1(net254009), .B2(n37749), .C1(net254201), .C2(n37746), 
        .A(n6577), .ZN(n6571) );
  OAI222_X1 U3481 ( .A1(n38022), .A2(n36050), .B1(n38370), .B2(n35538), .C1(
        n38195), .C2(n36562), .ZN(n6577) );
  AOI221_X1 U3482 ( .B1(net254297), .B2(n37725), .C1(net253881), .C2(n37722), 
        .A(n6586), .ZN(n6583) );
  OAI222_X1 U3483 ( .A1(n38271), .A2(n36051), .B1(n38088), .B2(n35539), .C1(
        n38444), .C2(n36563), .ZN(n6586) );
  AOI221_X1 U3484 ( .B1(net254010), .B2(n37749), .C1(net254202), .C2(n37746), 
        .A(n6535), .ZN(n6529) );
  OAI222_X1 U3485 ( .A1(n38022), .A2(n36052), .B1(n38370), .B2(n35540), .C1(
        n38195), .C2(n36564), .ZN(n6535) );
  AOI221_X1 U3486 ( .B1(net254298), .B2(n37725), .C1(net253882), .C2(n37722), 
        .A(n6544), .ZN(n6541) );
  OAI222_X1 U3487 ( .A1(n38271), .A2(n36053), .B1(n38088), .B2(n35541), .C1(
        n38444), .C2(n36565), .ZN(n6544) );
  AOI221_X1 U3488 ( .B1(net254011), .B2(n37750), .C1(net254203), .C2(n37747), 
        .A(n6365), .ZN(n6359) );
  OAI222_X1 U3489 ( .A1(n38022), .A2(n36054), .B1(n38370), .B2(n35542), .C1(
        n38196), .C2(n36566), .ZN(n6365) );
  AOI221_X1 U3490 ( .B1(net254299), .B2(n37726), .C1(net253883), .C2(n37723), 
        .A(n6444), .ZN(n6408) );
  OAI222_X1 U3491 ( .A1(n38271), .A2(n36055), .B1(n38088), .B2(n35543), .C1(
        n38445), .C2(n36567), .ZN(n6444) );
  AOI221_X1 U3492 ( .B1(net254012), .B2(n37750), .C1(net254204), .C2(n37747), 
        .A(n6323), .ZN(n6317) );
  OAI222_X1 U3493 ( .A1(n38022), .A2(n36056), .B1(n38370), .B2(n35544), .C1(
        n38196), .C2(n36568), .ZN(n6323) );
  AOI221_X1 U3494 ( .B1(net254300), .B2(n37726), .C1(net253884), .C2(n37723), 
        .A(n6332), .ZN(n6329) );
  OAI222_X1 U3495 ( .A1(n38271), .A2(n36057), .B1(n38088), .B2(n35545), .C1(
        n38445), .C2(n36569), .ZN(n6332) );
  AOI221_X1 U3496 ( .B1(net254013), .B2(n37750), .C1(net254205), .C2(n37747), 
        .A(n6281), .ZN(n6275) );
  OAI222_X1 U3497 ( .A1(n38022), .A2(n36058), .B1(n38370), .B2(n35546), .C1(
        n38196), .C2(n36570), .ZN(n6281) );
  AOI221_X1 U3498 ( .B1(net254301), .B2(n37726), .C1(net253885), .C2(n37723), 
        .A(n6290), .ZN(n6287) );
  OAI222_X1 U3499 ( .A1(n38271), .A2(n36059), .B1(n38088), .B2(n35547), .C1(
        n38445), .C2(n36571), .ZN(n6290) );
  AOI221_X1 U3500 ( .B1(net254014), .B2(n37750), .C1(net254206), .C2(n37747), 
        .A(n6239), .ZN(n6233) );
  OAI222_X1 U3501 ( .A1(n38022), .A2(n36060), .B1(n38370), .B2(n35548), .C1(
        n38196), .C2(n36572), .ZN(n6239) );
  AOI221_X1 U3502 ( .B1(net254302), .B2(n37726), .C1(net253886), .C2(n37723), 
        .A(n6248), .ZN(n6245) );
  OAI222_X1 U3503 ( .A1(n38271), .A2(n36061), .B1(n38088), .B2(n35549), .C1(
        n38445), .C2(n36573), .ZN(n6248) );
  AOI221_X1 U3504 ( .B1(net254015), .B2(n37750), .C1(net254207), .C2(n37747), 
        .A(n6197), .ZN(n6191) );
  OAI222_X1 U3505 ( .A1(n38022), .A2(n36062), .B1(n38370), .B2(n35550), .C1(
        n38196), .C2(n36574), .ZN(n6197) );
  AOI221_X1 U3506 ( .B1(net254303), .B2(n37726), .C1(net253887), .C2(n37723), 
        .A(n6206), .ZN(n6203) );
  OAI222_X1 U3507 ( .A1(n38271), .A2(n36063), .B1(n38088), .B2(n35551), .C1(
        n38445), .C2(n36575), .ZN(n6206) );
  AOI221_X1 U3508 ( .B1(net254016), .B2(n37750), .C1(net254208), .C2(n37747), 
        .A(n6155), .ZN(n6149) );
  OAI222_X1 U3509 ( .A1(n38022), .A2(n36064), .B1(n38370), .B2(n35552), .C1(
        n38196), .C2(n36576), .ZN(n6155) );
  AOI221_X1 U3510 ( .B1(net254304), .B2(n37726), .C1(net253888), .C2(n37723), 
        .A(n6164), .ZN(n6161) );
  OAI222_X1 U3511 ( .A1(n38271), .A2(n36065), .B1(n38088), .B2(n35553), .C1(
        n38445), .C2(n36577), .ZN(n6164) );
  AOI221_X1 U3512 ( .B1(net254017), .B2(n37750), .C1(net254209), .C2(n37747), 
        .A(n6113), .ZN(n6107) );
  OAI222_X1 U3513 ( .A1(n38022), .A2(n36066), .B1(n38370), .B2(n35554), .C1(
        n38196), .C2(n36578), .ZN(n6113) );
  AOI221_X1 U3514 ( .B1(net254305), .B2(n37726), .C1(net253889), .C2(n37723), 
        .A(n6122), .ZN(n6119) );
  OAI222_X1 U3515 ( .A1(n38271), .A2(n36067), .B1(n38088), .B2(n35555), .C1(
        n38445), .C2(n36579), .ZN(n6122) );
  AOI221_X1 U3516 ( .B1(net254018), .B2(n37750), .C1(net254210), .C2(n37747), 
        .A(n6071), .ZN(n6065) );
  OAI222_X1 U3517 ( .A1(n38022), .A2(n36068), .B1(n38370), .B2(n35556), .C1(
        n38196), .C2(n36580), .ZN(n6071) );
  AOI221_X1 U3518 ( .B1(net254306), .B2(n37726), .C1(net253890), .C2(n37723), 
        .A(n6080), .ZN(n6077) );
  OAI222_X1 U3519 ( .A1(n38271), .A2(n36069), .B1(n38088), .B2(n35557), .C1(
        n38445), .C2(n36581), .ZN(n6080) );
  AOI221_X1 U3520 ( .B1(net254019), .B2(n37750), .C1(net254211), .C2(n37747), 
        .A(n6029), .ZN(n6023) );
  OAI222_X1 U3521 ( .A1(n38022), .A2(n36070), .B1(n38370), .B2(n35558), .C1(
        n38196), .C2(n36582), .ZN(n6029) );
  AOI221_X1 U3522 ( .B1(net254307), .B2(n37726), .C1(net253891), .C2(n37723), 
        .A(n6038), .ZN(n6035) );
  OAI222_X1 U3523 ( .A1(n38271), .A2(n36071), .B1(n38088), .B2(n35559), .C1(
        n38445), .C2(n36583), .ZN(n6038) );
  AOI221_X1 U3524 ( .B1(net254020), .B2(n37750), .C1(net254212), .C2(n37747), 
        .A(n5987), .ZN(n5981) );
  OAI222_X1 U3525 ( .A1(n38021), .A2(n36072), .B1(n38369), .B2(n35560), .C1(
        n38196), .C2(n36584), .ZN(n5987) );
  AOI221_X1 U3526 ( .B1(net254308), .B2(n37726), .C1(net253892), .C2(n37723), 
        .A(n5996), .ZN(n5993) );
  OAI222_X1 U3527 ( .A1(n38270), .A2(n36073), .B1(n38087), .B2(n35561), .C1(
        n38445), .C2(n36585), .ZN(n5996) );
  AOI221_X1 U3528 ( .B1(net254021), .B2(n37750), .C1(net254213), .C2(n37747), 
        .A(n5945), .ZN(n5939) );
  OAI222_X1 U3529 ( .A1(n38021), .A2(n36074), .B1(n38369), .B2(n35562), .C1(
        n38196), .C2(n36586), .ZN(n5945) );
  AOI221_X1 U3530 ( .B1(net254309), .B2(n37726), .C1(net253893), .C2(n37723), 
        .A(n5954), .ZN(n5951) );
  OAI222_X1 U3531 ( .A1(n38270), .A2(n36075), .B1(n38087), .B2(n35563), .C1(
        n38445), .C2(n36587), .ZN(n5954) );
  AOI221_X1 U3532 ( .B1(net254022), .B2(n37750), .C1(net254214), .C2(n37747), 
        .A(n5903), .ZN(n5897) );
  OAI222_X1 U3533 ( .A1(n38021), .A2(n36076), .B1(n38369), .B2(n35564), .C1(
        n38196), .C2(n36588), .ZN(n5903) );
  AOI221_X1 U3534 ( .B1(net254310), .B2(n37726), .C1(net253894), .C2(n37723), 
        .A(n5912), .ZN(n5909) );
  OAI222_X1 U3535 ( .A1(n38270), .A2(n36077), .B1(n38087), .B2(n35565), .C1(
        n38445), .C2(n36589), .ZN(n5912) );
  AOI221_X1 U3536 ( .B1(net253935), .B2(n37743), .C1(net254127), .C2(n37740), 
        .A(n9617), .ZN(n9608) );
  OAI222_X1 U3537 ( .A1(n37969), .A2(n36078), .B1(n38317), .B2(n35566), .C1(
        n38141), .C2(n36590), .ZN(n9617) );
  AOI221_X1 U3538 ( .B1(net254223), .B2(n37719), .C1(net253807), .C2(n37716), 
        .A(n9627), .ZN(n9621) );
  OAI222_X1 U3539 ( .A1(n38218), .A2(n36079), .B1(n38035), .B2(n35567), .C1(
        n38390), .C2(n36591), .ZN(n9627) );
  AOI221_X1 U3540 ( .B1(net253936), .B2(n37743), .C1(net254128), .C2(n37740), 
        .A(n9549), .ZN(n9540) );
  OAI222_X1 U3541 ( .A1(n37969), .A2(n36080), .B1(n38317), .B2(n35568), .C1(
        n38141), .C2(n36592), .ZN(n9549) );
  AOI221_X1 U3542 ( .B1(net254224), .B2(n37719), .C1(net253808), .C2(n37716), 
        .A(n9557), .ZN(n9552) );
  OAI222_X1 U3543 ( .A1(n38218), .A2(n36081), .B1(n38035), .B2(n35569), .C1(
        n38390), .C2(n36593), .ZN(n9557) );
  AOI221_X1 U3544 ( .B1(net253937), .B2(n37743), .C1(net254129), .C2(n37740), 
        .A(n9507), .ZN(n9498) );
  OAI222_X1 U3545 ( .A1(n37969), .A2(n36082), .B1(n38317), .B2(n35570), .C1(
        n38141), .C2(n36594), .ZN(n9507) );
  AOI221_X1 U3546 ( .B1(net254225), .B2(n37719), .C1(net253809), .C2(n37716), 
        .A(n9515), .ZN(n9510) );
  OAI222_X1 U3547 ( .A1(n38218), .A2(n36083), .B1(n38035), .B2(n35571), .C1(
        n38390), .C2(n36595), .ZN(n9515) );
  AOI221_X1 U3548 ( .B1(net253938), .B2(n37743), .C1(net254130), .C2(n37740), 
        .A(n9465), .ZN(n9456) );
  OAI222_X1 U3549 ( .A1(n37969), .A2(n36084), .B1(n38317), .B2(n35572), .C1(
        n38141), .C2(n36596), .ZN(n9465) );
  AOI221_X1 U3550 ( .B1(net254226), .B2(n37719), .C1(net253810), .C2(n37716), 
        .A(n9473), .ZN(n9468) );
  OAI222_X1 U3551 ( .A1(n38218), .A2(n36085), .B1(n38035), .B2(n35573), .C1(
        n38390), .C2(n36597), .ZN(n9473) );
  AOI221_X1 U3552 ( .B1(net253939), .B2(n37743), .C1(net254131), .C2(n37740), 
        .A(n9423), .ZN(n9414) );
  OAI222_X1 U3553 ( .A1(n37969), .A2(n36086), .B1(n38317), .B2(n35574), .C1(
        n38141), .C2(n36598), .ZN(n9423) );
  AOI221_X1 U3554 ( .B1(net254227), .B2(n37719), .C1(net253811), .C2(n37716), 
        .A(n9431), .ZN(n9426) );
  OAI222_X1 U3555 ( .A1(n38218), .A2(n36087), .B1(n38035), .B2(n35575), .C1(
        n38390), .C2(n36599), .ZN(n9431) );
  AOI221_X1 U3556 ( .B1(net253940), .B2(n37743), .C1(net254132), .C2(n37740), 
        .A(n9381), .ZN(n9372) );
  OAI222_X1 U3557 ( .A1(n37969), .A2(n36088), .B1(n38317), .B2(n35576), .C1(
        n38141), .C2(n36600), .ZN(n9381) );
  AOI221_X1 U3558 ( .B1(net254228), .B2(n37719), .C1(net253812), .C2(n37716), 
        .A(n9389), .ZN(n9384) );
  OAI222_X1 U3559 ( .A1(n38218), .A2(n36089), .B1(n38035), .B2(n35577), .C1(
        n38390), .C2(n36601), .ZN(n9389) );
  AOI221_X1 U3560 ( .B1(net253941), .B2(n37743), .C1(net254133), .C2(n37740), 
        .A(n9339), .ZN(n9330) );
  OAI222_X1 U3561 ( .A1(n37969), .A2(n36090), .B1(n38317), .B2(n35578), .C1(
        n38141), .C2(n36602), .ZN(n9339) );
  AOI221_X1 U3562 ( .B1(net254229), .B2(n37719), .C1(net253813), .C2(n37716), 
        .A(n9347), .ZN(n9342) );
  OAI222_X1 U3563 ( .A1(n38218), .A2(n36091), .B1(n38035), .B2(n35579), .C1(
        n38390), .C2(n36603), .ZN(n9347) );
  AOI221_X1 U3564 ( .B1(net253942), .B2(n37743), .C1(net254134), .C2(n37740), 
        .A(n9297), .ZN(n9288) );
  OAI222_X1 U3565 ( .A1(n37969), .A2(n36092), .B1(n38317), .B2(n35580), .C1(
        n38141), .C2(n36604), .ZN(n9297) );
  AOI221_X1 U3566 ( .B1(net254230), .B2(n37719), .C1(net253814), .C2(n37716), 
        .A(n9305), .ZN(n9300) );
  OAI222_X1 U3567 ( .A1(n38218), .A2(n36093), .B1(n38035), .B2(n35581), .C1(
        n38390), .C2(n36605), .ZN(n9305) );
  AOI221_X1 U3568 ( .B1(net253943), .B2(n37743), .C1(net254135), .C2(n37740), 
        .A(n6663), .ZN(n6654) );
  OAI222_X1 U3569 ( .A1(n37969), .A2(n36094), .B1(n38317), .B2(n35582), .C1(
        n38141), .C2(n36606), .ZN(n6663) );
  AOI221_X1 U3570 ( .B1(net254231), .B2(n37719), .C1(net253815), .C2(n37716), 
        .A(n6671), .ZN(n6666) );
  OAI222_X1 U3571 ( .A1(n38218), .A2(n36095), .B1(n38035), .B2(n35583), .C1(
        n38390), .C2(n36607), .ZN(n6671) );
  AOI221_X1 U3572 ( .B1(net253944), .B2(n37743), .C1(net254136), .C2(n37740), 
        .A(n6621), .ZN(n6612) );
  OAI222_X1 U3573 ( .A1(n37968), .A2(n36096), .B1(n38316), .B2(n35584), .C1(
        n38141), .C2(n36608), .ZN(n6621) );
  AOI221_X1 U3574 ( .B1(net254232), .B2(n37719), .C1(net253816), .C2(n37716), 
        .A(n6629), .ZN(n6624) );
  OAI222_X1 U3575 ( .A1(n38217), .A2(n36097), .B1(n38034), .B2(n35585), .C1(
        n38390), .C2(n36609), .ZN(n6629) );
  AOI221_X1 U3576 ( .B1(net253945), .B2(n37743), .C1(net254137), .C2(n37740), 
        .A(n6579), .ZN(n6570) );
  OAI222_X1 U3577 ( .A1(n37968), .A2(n36098), .B1(n38316), .B2(n35586), .C1(
        n38141), .C2(n36610), .ZN(n6579) );
  AOI221_X1 U3578 ( .B1(net254233), .B2(n37719), .C1(net253817), .C2(n37716), 
        .A(n6587), .ZN(n6582) );
  OAI222_X1 U3579 ( .A1(n38217), .A2(n36099), .B1(n38034), .B2(n35587), .C1(
        n38390), .C2(n36611), .ZN(n6587) );
  AOI221_X1 U3580 ( .B1(net253946), .B2(n37743), .C1(net254138), .C2(n37740), 
        .A(n6537), .ZN(n6528) );
  OAI222_X1 U3581 ( .A1(n37968), .A2(n36100), .B1(n38316), .B2(n35588), .C1(
        n38141), .C2(n36612), .ZN(n6537) );
  AOI221_X1 U3582 ( .B1(net254234), .B2(n37719), .C1(net253818), .C2(n37716), 
        .A(n6545), .ZN(n6540) );
  OAI222_X1 U3583 ( .A1(n38217), .A2(n36101), .B1(n38034), .B2(n35589), .C1(
        n38390), .C2(n36613), .ZN(n6545) );
  AOI221_X1 U3584 ( .B1(net253947), .B2(n37744), .C1(net254139), .C2(n37741), 
        .A(n6367), .ZN(n6358) );
  OAI222_X1 U3585 ( .A1(n37968), .A2(n36102), .B1(n38316), .B2(n35590), .C1(
        n38142), .C2(n36614), .ZN(n6367) );
  AOI221_X1 U3586 ( .B1(net254235), .B2(n37720), .C1(net253819), .C2(n37717), 
        .A(n6446), .ZN(n6406) );
  OAI222_X1 U3587 ( .A1(n38217), .A2(n36103), .B1(n38034), .B2(n35591), .C1(
        n38391), .C2(n36615), .ZN(n6446) );
  AOI221_X1 U3588 ( .B1(net253948), .B2(n37744), .C1(net254140), .C2(n37741), 
        .A(n6325), .ZN(n6316) );
  OAI222_X1 U3589 ( .A1(n37968), .A2(n36104), .B1(n38316), .B2(n35592), .C1(
        n38142), .C2(n36616), .ZN(n6325) );
  AOI221_X1 U3590 ( .B1(net254236), .B2(n37720), .C1(net253820), .C2(n37717), 
        .A(n6333), .ZN(n6328) );
  OAI222_X1 U3591 ( .A1(n38217), .A2(n36105), .B1(n38034), .B2(n35593), .C1(
        n38391), .C2(n36617), .ZN(n6333) );
  AOI221_X1 U3592 ( .B1(net253949), .B2(n37744), .C1(net254141), .C2(n37741), 
        .A(n6283), .ZN(n6274) );
  OAI222_X1 U3593 ( .A1(n37968), .A2(n36106), .B1(n38316), .B2(n35594), .C1(
        n38142), .C2(n36618), .ZN(n6283) );
  AOI221_X1 U3594 ( .B1(net254237), .B2(n37720), .C1(net253821), .C2(n37717), 
        .A(n6291), .ZN(n6286) );
  OAI222_X1 U3595 ( .A1(n38217), .A2(n36107), .B1(n38034), .B2(n35595), .C1(
        n38391), .C2(n36619), .ZN(n6291) );
  AOI221_X1 U3596 ( .B1(net253950), .B2(n37744), .C1(net254142), .C2(n37741), 
        .A(n6241), .ZN(n6232) );
  OAI222_X1 U3597 ( .A1(n37968), .A2(n36108), .B1(n38316), .B2(n35596), .C1(
        n38142), .C2(n36620), .ZN(n6241) );
  AOI221_X1 U3598 ( .B1(net254238), .B2(n37720), .C1(net253822), .C2(n37717), 
        .A(n6249), .ZN(n6244) );
  OAI222_X1 U3599 ( .A1(n38217), .A2(n36109), .B1(n38034), .B2(n35597), .C1(
        n38391), .C2(n36621), .ZN(n6249) );
  AOI221_X1 U3600 ( .B1(net253951), .B2(n37744), .C1(net254143), .C2(n37741), 
        .A(n6199), .ZN(n6190) );
  OAI222_X1 U3601 ( .A1(n37968), .A2(n36110), .B1(n38316), .B2(n35598), .C1(
        n38142), .C2(n36622), .ZN(n6199) );
  AOI221_X1 U3602 ( .B1(net254239), .B2(n37720), .C1(net253823), .C2(n37717), 
        .A(n6207), .ZN(n6202) );
  OAI222_X1 U3603 ( .A1(n38217), .A2(n36111), .B1(n38034), .B2(n35599), .C1(
        n38391), .C2(n36623), .ZN(n6207) );
  AOI221_X1 U3604 ( .B1(net253952), .B2(n37744), .C1(net254144), .C2(n37741), 
        .A(n6157), .ZN(n6148) );
  OAI222_X1 U3605 ( .A1(n37968), .A2(n36112), .B1(n38316), .B2(n35600), .C1(
        n38142), .C2(n36624), .ZN(n6157) );
  AOI221_X1 U3606 ( .B1(net254240), .B2(n37720), .C1(net253824), .C2(n37717), 
        .A(n6165), .ZN(n6160) );
  OAI222_X1 U3607 ( .A1(n38217), .A2(n36113), .B1(n38034), .B2(n35601), .C1(
        n38391), .C2(n36625), .ZN(n6165) );
  AOI221_X1 U3608 ( .B1(net253953), .B2(n37744), .C1(net254145), .C2(n37741), 
        .A(n6115), .ZN(n6106) );
  OAI222_X1 U3609 ( .A1(n37968), .A2(n36114), .B1(n38316), .B2(n35602), .C1(
        n38142), .C2(n36626), .ZN(n6115) );
  AOI221_X1 U3610 ( .B1(net254241), .B2(n37720), .C1(net253825), .C2(n37717), 
        .A(n6123), .ZN(n6118) );
  OAI222_X1 U3611 ( .A1(n38217), .A2(n36115), .B1(n38034), .B2(n35603), .C1(
        n38391), .C2(n36627), .ZN(n6123) );
  AOI221_X1 U3612 ( .B1(net253954), .B2(n37744), .C1(net254146), .C2(n37741), 
        .A(n6073), .ZN(n6064) );
  OAI222_X1 U3613 ( .A1(n37968), .A2(n36116), .B1(n38316), .B2(n35604), .C1(
        n38142), .C2(n36628), .ZN(n6073) );
  AOI221_X1 U3614 ( .B1(net254242), .B2(n37720), .C1(net253826), .C2(n37717), 
        .A(n6081), .ZN(n6076) );
  OAI222_X1 U3615 ( .A1(n38217), .A2(n36117), .B1(n38034), .B2(n35605), .C1(
        n38391), .C2(n36629), .ZN(n6081) );
  AOI221_X1 U3616 ( .B1(net253955), .B2(n37744), .C1(net254147), .C2(n37741), 
        .A(n6031), .ZN(n6022) );
  OAI222_X1 U3617 ( .A1(n37968), .A2(n36118), .B1(n38316), .B2(n35606), .C1(
        n38142), .C2(n36630), .ZN(n6031) );
  AOI221_X1 U3618 ( .B1(net254243), .B2(n37720), .C1(net253827), .C2(n37717), 
        .A(n6039), .ZN(n6034) );
  OAI222_X1 U3619 ( .A1(n38217), .A2(n36119), .B1(n38034), .B2(n35607), .C1(
        n38391), .C2(n36631), .ZN(n6039) );
  AOI221_X1 U3620 ( .B1(net253956), .B2(n37744), .C1(net254148), .C2(n37741), 
        .A(n5989), .ZN(n5980) );
  OAI222_X1 U3621 ( .A1(n37967), .A2(n36120), .B1(n38315), .B2(n35608), .C1(
        n38142), .C2(n36632), .ZN(n5989) );
  AOI221_X1 U3622 ( .B1(net254244), .B2(n37720), .C1(net253828), .C2(n37717), 
        .A(n5997), .ZN(n5992) );
  OAI222_X1 U3623 ( .A1(n38216), .A2(n36121), .B1(n38033), .B2(n35609), .C1(
        n38391), .C2(n36633), .ZN(n5997) );
  AOI221_X1 U3624 ( .B1(net253957), .B2(n37744), .C1(net254149), .C2(n37741), 
        .A(n5947), .ZN(n5938) );
  OAI222_X1 U3625 ( .A1(n37967), .A2(n36122), .B1(n38315), .B2(n35610), .C1(
        n38142), .C2(n36634), .ZN(n5947) );
  AOI221_X1 U3626 ( .B1(net254245), .B2(n37720), .C1(net253829), .C2(n37717), 
        .A(n5955), .ZN(n5950) );
  OAI222_X1 U3627 ( .A1(n38216), .A2(n36123), .B1(n38033), .B2(n35611), .C1(
        n38391), .C2(n36635), .ZN(n5955) );
  AOI221_X1 U3628 ( .B1(net253958), .B2(n37744), .C1(net254150), .C2(n37741), 
        .A(n5905), .ZN(n5896) );
  OAI222_X1 U3629 ( .A1(n37967), .A2(n36124), .B1(n38315), .B2(n35612), .C1(
        n38142), .C2(n36636), .ZN(n5905) );
  AOI221_X1 U3630 ( .B1(net254246), .B2(n37720), .C1(net253830), .C2(n37717), 
        .A(n5913), .ZN(n5908) );
  OAI222_X1 U3631 ( .A1(n38216), .A2(n36125), .B1(n38033), .B2(n35613), .C1(
        n38391), .C2(n36637), .ZN(n5913) );
  AOI221_X1 U3632 ( .B1(net254159), .B2(n37737), .C1(net253743), .C2(n37734), 
        .A(n9618), .ZN(n9607) );
  OAI222_X1 U3633 ( .A1(n38164), .A2(n36126), .B1(n37981), .B2(n35614), .C1(
        n38336), .C2(n36638), .ZN(n9618) );
  AOI221_X1 U3634 ( .B1(net253839), .B2(n37713), .C1(net254031), .C2(n37710), 
        .A(n9628), .ZN(n9620) );
  OAI222_X1 U3635 ( .A1(n38413), .A2(n36127), .B1(n38230), .B2(n35615), .C1(
        n38054), .C2(n36639), .ZN(n9628) );
  AOI221_X1 U3636 ( .B1(net254160), .B2(n37737), .C1(net253744), .C2(n37734), 
        .A(n9550), .ZN(n9539) );
  OAI222_X1 U3637 ( .A1(n38164), .A2(n36128), .B1(n37981), .B2(n35616), .C1(
        n38336), .C2(n36640), .ZN(n9550) );
  AOI221_X1 U3638 ( .B1(net253840), .B2(n37713), .C1(net254032), .C2(n37710), 
        .A(n9558), .ZN(n9551) );
  OAI222_X1 U3639 ( .A1(n38413), .A2(n36129), .B1(n38230), .B2(n35617), .C1(
        n38054), .C2(n36641), .ZN(n9558) );
  AOI221_X1 U3640 ( .B1(net254161), .B2(n37737), .C1(net253745), .C2(n37734), 
        .A(n9508), .ZN(n9497) );
  OAI222_X1 U3641 ( .A1(n38164), .A2(n36130), .B1(n37981), .B2(n35618), .C1(
        n38336), .C2(n36642), .ZN(n9508) );
  AOI221_X1 U3642 ( .B1(net253841), .B2(n37713), .C1(net254033), .C2(n37710), 
        .A(n9516), .ZN(n9509) );
  OAI222_X1 U3643 ( .A1(n38413), .A2(n36131), .B1(n38230), .B2(n35619), .C1(
        n38054), .C2(n36643), .ZN(n9516) );
  AOI221_X1 U3644 ( .B1(net254162), .B2(n37737), .C1(net253746), .C2(n37734), 
        .A(n9466), .ZN(n9455) );
  OAI222_X1 U3645 ( .A1(n38164), .A2(n36132), .B1(n37981), .B2(n35620), .C1(
        n38336), .C2(n36644), .ZN(n9466) );
  AOI221_X1 U3646 ( .B1(net253842), .B2(n37713), .C1(net254034), .C2(n37710), 
        .A(n9474), .ZN(n9467) );
  OAI222_X1 U3647 ( .A1(n38413), .A2(n36133), .B1(n38230), .B2(n35621), .C1(
        n38054), .C2(n36645), .ZN(n9474) );
  AOI221_X1 U3648 ( .B1(net254163), .B2(n37737), .C1(net253747), .C2(n37734), 
        .A(n9424), .ZN(n9413) );
  OAI222_X1 U3649 ( .A1(n38164), .A2(n36134), .B1(n37981), .B2(n35622), .C1(
        n38336), .C2(n36646), .ZN(n9424) );
  AOI221_X1 U3650 ( .B1(net253843), .B2(n37713), .C1(net254035), .C2(n37710), 
        .A(n9432), .ZN(n9425) );
  OAI222_X1 U3651 ( .A1(n38413), .A2(n36135), .B1(n38230), .B2(n35623), .C1(
        n38054), .C2(n36647), .ZN(n9432) );
  AOI221_X1 U3652 ( .B1(net254164), .B2(n37737), .C1(net253748), .C2(n37734), 
        .A(n9382), .ZN(n9371) );
  OAI222_X1 U3653 ( .A1(n38164), .A2(n36136), .B1(n37981), .B2(n35624), .C1(
        n38336), .C2(n36648), .ZN(n9382) );
  AOI221_X1 U3654 ( .B1(net253844), .B2(n37713), .C1(net254036), .C2(n37710), 
        .A(n9390), .ZN(n9383) );
  OAI222_X1 U3655 ( .A1(n38413), .A2(n36137), .B1(n38230), .B2(n35625), .C1(
        n38054), .C2(n36649), .ZN(n9390) );
  AOI221_X1 U3656 ( .B1(net254165), .B2(n37737), .C1(net253749), .C2(n37734), 
        .A(n9340), .ZN(n9329) );
  OAI222_X1 U3657 ( .A1(n38164), .A2(n36138), .B1(n37981), .B2(n35626), .C1(
        n38336), .C2(n36650), .ZN(n9340) );
  AOI221_X1 U3658 ( .B1(net253845), .B2(n37713), .C1(net254037), .C2(n37710), 
        .A(n9348), .ZN(n9341) );
  OAI222_X1 U3659 ( .A1(n38413), .A2(n36139), .B1(n38230), .B2(n35627), .C1(
        n38054), .C2(n36651), .ZN(n9348) );
  AOI221_X1 U3660 ( .B1(net254166), .B2(n37737), .C1(net253750), .C2(n37734), 
        .A(n9298), .ZN(n9287) );
  OAI222_X1 U3661 ( .A1(n38164), .A2(n36140), .B1(n37981), .B2(n35628), .C1(
        n38336), .C2(n36652), .ZN(n9298) );
  AOI221_X1 U3662 ( .B1(net253846), .B2(n37713), .C1(net254038), .C2(n37710), 
        .A(n9306), .ZN(n9299) );
  OAI222_X1 U3663 ( .A1(n38413), .A2(n36141), .B1(n38230), .B2(n35629), .C1(
        n38054), .C2(n36653), .ZN(n9306) );
  AOI221_X1 U3664 ( .B1(net254167), .B2(n37737), .C1(net253751), .C2(n37734), 
        .A(n6664), .ZN(n6653) );
  OAI222_X1 U3665 ( .A1(n38164), .A2(n36142), .B1(n37981), .B2(n35630), .C1(
        n38336), .C2(n36654), .ZN(n6664) );
  AOI221_X1 U3666 ( .B1(net253847), .B2(n37713), .C1(net254039), .C2(n37710), 
        .A(n6672), .ZN(n6665) );
  OAI222_X1 U3667 ( .A1(n38413), .A2(n36143), .B1(n38230), .B2(n35631), .C1(
        n38054), .C2(n36655), .ZN(n6672) );
  AOI221_X1 U3668 ( .B1(net254168), .B2(n37737), .C1(net253752), .C2(n37734), 
        .A(n6622), .ZN(n6611) );
  OAI222_X1 U3669 ( .A1(n38163), .A2(n36144), .B1(n37980), .B2(n35632), .C1(
        n38336), .C2(n36656), .ZN(n6622) );
  AOI221_X1 U3670 ( .B1(net253848), .B2(n37713), .C1(net254040), .C2(n37710), 
        .A(n6630), .ZN(n6623) );
  OAI222_X1 U3671 ( .A1(n38412), .A2(n36145), .B1(n38229), .B2(n35633), .C1(
        n38054), .C2(n36657), .ZN(n6630) );
  AOI221_X1 U3672 ( .B1(net254169), .B2(n37737), .C1(net253753), .C2(n37734), 
        .A(n6580), .ZN(n6569) );
  OAI222_X1 U3673 ( .A1(n38163), .A2(n36146), .B1(n37980), .B2(n35634), .C1(
        n38336), .C2(n36658), .ZN(n6580) );
  AOI221_X1 U3674 ( .B1(net253849), .B2(n37713), .C1(net254041), .C2(n37710), 
        .A(n6588), .ZN(n6581) );
  OAI222_X1 U3675 ( .A1(n38412), .A2(n36147), .B1(n38229), .B2(n35635), .C1(
        n38054), .C2(n36659), .ZN(n6588) );
  AOI221_X1 U3676 ( .B1(net254170), .B2(n37737), .C1(net253754), .C2(n37734), 
        .A(n6538), .ZN(n6527) );
  OAI222_X1 U3677 ( .A1(n38163), .A2(n36148), .B1(n37980), .B2(n35636), .C1(
        n38336), .C2(n36660), .ZN(n6538) );
  AOI221_X1 U3678 ( .B1(net253850), .B2(n37713), .C1(net254042), .C2(n37710), 
        .A(n6546), .ZN(n6539) );
  OAI222_X1 U3679 ( .A1(n38412), .A2(n36149), .B1(n38229), .B2(n35637), .C1(
        n38054), .C2(n36661), .ZN(n6546) );
  AOI221_X1 U3680 ( .B1(net254171), .B2(n37738), .C1(net253755), .C2(n37735), 
        .A(n6371), .ZN(n6357) );
  OAI222_X1 U3681 ( .A1(n38163), .A2(n36150), .B1(n37980), .B2(n35638), .C1(
        n38337), .C2(n36662), .ZN(n6371) );
  AOI221_X1 U3682 ( .B1(net253851), .B2(n37714), .C1(net254043), .C2(n37711), 
        .A(n6447), .ZN(n6373) );
  OAI222_X1 U3683 ( .A1(n38412), .A2(n36151), .B1(n38229), .B2(n35639), .C1(
        n38055), .C2(n36663), .ZN(n6447) );
  AOI221_X1 U3684 ( .B1(net254172), .B2(n37738), .C1(net253756), .C2(n37735), 
        .A(n6326), .ZN(n6315) );
  OAI222_X1 U3685 ( .A1(n38163), .A2(n36152), .B1(n37980), .B2(n35640), .C1(
        n38337), .C2(n36664), .ZN(n6326) );
  AOI221_X1 U3686 ( .B1(net253852), .B2(n37714), .C1(net254044), .C2(n37711), 
        .A(n6334), .ZN(n6327) );
  OAI222_X1 U3687 ( .A1(n38412), .A2(n36153), .B1(n38229), .B2(n35641), .C1(
        n38055), .C2(n36665), .ZN(n6334) );
  AOI221_X1 U3688 ( .B1(net254173), .B2(n37738), .C1(net253757), .C2(n37735), 
        .A(n6284), .ZN(n6273) );
  OAI222_X1 U3689 ( .A1(n38163), .A2(n36154), .B1(n37980), .B2(n35642), .C1(
        n38337), .C2(n36666), .ZN(n6284) );
  AOI221_X1 U3690 ( .B1(net253853), .B2(n37714), .C1(net254045), .C2(n37711), 
        .A(n6292), .ZN(n6285) );
  OAI222_X1 U3691 ( .A1(n38412), .A2(n36155), .B1(n38229), .B2(n35643), .C1(
        n38055), .C2(n36667), .ZN(n6292) );
  AOI221_X1 U3692 ( .B1(net254174), .B2(n37738), .C1(net253758), .C2(n37735), 
        .A(n6242), .ZN(n6231) );
  OAI222_X1 U3693 ( .A1(n38163), .A2(n36156), .B1(n37980), .B2(n35644), .C1(
        n38337), .C2(n36668), .ZN(n6242) );
  AOI221_X1 U3694 ( .B1(net253854), .B2(n37714), .C1(net254046), .C2(n37711), 
        .A(n6250), .ZN(n6243) );
  OAI222_X1 U3695 ( .A1(n38412), .A2(n36157), .B1(n38229), .B2(n35645), .C1(
        n38055), .C2(n36669), .ZN(n6250) );
  AOI221_X1 U3696 ( .B1(net254175), .B2(n37738), .C1(net253759), .C2(n37735), 
        .A(n6200), .ZN(n6189) );
  OAI222_X1 U3697 ( .A1(n38163), .A2(n36158), .B1(n37980), .B2(n35646), .C1(
        n38337), .C2(n36670), .ZN(n6200) );
  AOI221_X1 U3698 ( .B1(net253855), .B2(n37714), .C1(net254047), .C2(n37711), 
        .A(n6208), .ZN(n6201) );
  OAI222_X1 U3699 ( .A1(n38412), .A2(n36159), .B1(n38229), .B2(n35647), .C1(
        n38055), .C2(n36671), .ZN(n6208) );
  AOI221_X1 U3700 ( .B1(net254176), .B2(n37738), .C1(net253760), .C2(n37735), 
        .A(n6158), .ZN(n6147) );
  OAI222_X1 U3701 ( .A1(n38163), .A2(n36160), .B1(n37980), .B2(n35648), .C1(
        n38337), .C2(n36672), .ZN(n6158) );
  AOI221_X1 U3702 ( .B1(net253856), .B2(n37714), .C1(net254048), .C2(n37711), 
        .A(n6166), .ZN(n6159) );
  OAI222_X1 U3703 ( .A1(n38412), .A2(n36161), .B1(n38229), .B2(n35649), .C1(
        n38055), .C2(n36673), .ZN(n6166) );
  AOI221_X1 U3704 ( .B1(net254177), .B2(n37738), .C1(net253761), .C2(n37735), 
        .A(n6116), .ZN(n6105) );
  OAI222_X1 U3705 ( .A1(n38163), .A2(n36162), .B1(n37980), .B2(n35650), .C1(
        n38337), .C2(n36674), .ZN(n6116) );
  AOI221_X1 U3706 ( .B1(net253857), .B2(n37714), .C1(net254049), .C2(n37711), 
        .A(n6124), .ZN(n6117) );
  OAI222_X1 U3707 ( .A1(n38412), .A2(n36163), .B1(n38229), .B2(n35651), .C1(
        n38055), .C2(n36675), .ZN(n6124) );
  AOI221_X1 U3708 ( .B1(net254178), .B2(n37738), .C1(net253762), .C2(n37735), 
        .A(n6074), .ZN(n6063) );
  OAI222_X1 U3709 ( .A1(n38163), .A2(n36164), .B1(n37980), .B2(n35652), .C1(
        n38337), .C2(n36676), .ZN(n6074) );
  AOI221_X1 U3710 ( .B1(net253858), .B2(n37714), .C1(net254050), .C2(n37711), 
        .A(n6082), .ZN(n6075) );
  OAI222_X1 U3711 ( .A1(n38412), .A2(n36165), .B1(n38229), .B2(n35653), .C1(
        n38055), .C2(n36677), .ZN(n6082) );
  AOI221_X1 U3712 ( .B1(net254179), .B2(n37738), .C1(net253763), .C2(n37735), 
        .A(n6032), .ZN(n6021) );
  OAI222_X1 U3713 ( .A1(n38163), .A2(n36166), .B1(n37980), .B2(n35654), .C1(
        n38337), .C2(n36678), .ZN(n6032) );
  AOI221_X1 U3714 ( .B1(net253859), .B2(n37714), .C1(net254051), .C2(n37711), 
        .A(n6040), .ZN(n6033) );
  OAI222_X1 U3715 ( .A1(n38412), .A2(n36167), .B1(n38229), .B2(n35655), .C1(
        n38055), .C2(n36679), .ZN(n6040) );
  AOI221_X1 U3716 ( .B1(net254180), .B2(n37738), .C1(net253764), .C2(n37735), 
        .A(n5990), .ZN(n5979) );
  OAI222_X1 U3717 ( .A1(n38162), .A2(n36168), .B1(n37979), .B2(n35656), .C1(
        n38337), .C2(n36680), .ZN(n5990) );
  AOI221_X1 U3718 ( .B1(net253860), .B2(n37714), .C1(net254052), .C2(n37711), 
        .A(n5998), .ZN(n5991) );
  OAI222_X1 U3719 ( .A1(n38411), .A2(n36169), .B1(n38228), .B2(n35657), .C1(
        n38055), .C2(n36681), .ZN(n5998) );
  AOI221_X1 U3720 ( .B1(net254181), .B2(n37738), .C1(net253765), .C2(n37735), 
        .A(n5948), .ZN(n5937) );
  OAI222_X1 U3721 ( .A1(n38162), .A2(n36170), .B1(n37979), .B2(n35658), .C1(
        n38337), .C2(n36682), .ZN(n5948) );
  AOI221_X1 U3722 ( .B1(net253861), .B2(n37714), .C1(net254053), .C2(n37711), 
        .A(n5956), .ZN(n5949) );
  OAI222_X1 U3723 ( .A1(n38411), .A2(n36171), .B1(n38228), .B2(n35659), .C1(
        n38055), .C2(n36683), .ZN(n5956) );
  AOI221_X1 U3724 ( .B1(net254182), .B2(n37738), .C1(net253766), .C2(n37735), 
        .A(n5906), .ZN(n5895) );
  OAI222_X1 U3725 ( .A1(n38162), .A2(n36172), .B1(n37979), .B2(n35660), .C1(
        n38337), .C2(n36684), .ZN(n5906) );
  AOI221_X1 U3726 ( .B1(net253862), .B2(n37714), .C1(net254054), .C2(n37711), 
        .A(n5914), .ZN(n5907) );
  OAI222_X1 U3727 ( .A1(n38411), .A2(n36173), .B1(n38228), .B2(n35661), .C1(
        n38055), .C2(n36685), .ZN(n5914) );
  OR3_X1 U3728 ( .A1(Addr[4]), .A2(Addr[5]), .A3(n2812), .ZN(n5016) );
  OAI22_X1 U3729 ( .A1(n38499), .A2(n37582), .B1(n38684), .B2(n38498), .ZN(
        n8755) );
  OAI22_X1 U3730 ( .A1(n38499), .A2(n37583), .B1(n38691), .B2(n38498), .ZN(
        n8756) );
  OAI22_X1 U3731 ( .A1(n38499), .A2(n37584), .B1(n38698), .B2(n38498), .ZN(
        n8757) );
  OAI22_X1 U3732 ( .A1(n38499), .A2(n37585), .B1(n38705), .B2(n38498), .ZN(
        n8758) );
  OAI22_X1 U3733 ( .A1(n38499), .A2(n37586), .B1(n38712), .B2(n38498), .ZN(
        n8759) );
  OAI22_X1 U3734 ( .A1(n38500), .A2(n37587), .B1(n38719), .B2(n38498), .ZN(
        n8760) );
  OAI22_X1 U3735 ( .A1(n38500), .A2(n37588), .B1(n38726), .B2(n38498), .ZN(
        n8761) );
  OAI22_X1 U3736 ( .A1(n38500), .A2(n37589), .B1(n38733), .B2(n38498), .ZN(
        n8762) );
  OAI22_X1 U3737 ( .A1(n38500), .A2(n37590), .B1(n38740), .B2(n38498), .ZN(
        n8763) );
  OAI22_X1 U3738 ( .A1(n38500), .A2(n37591), .B1(n38747), .B2(n38498), .ZN(
        n8764) );
  OAI22_X1 U3739 ( .A1(n38501), .A2(n37592), .B1(n38754), .B2(n38498), .ZN(
        n8765) );
  OAI22_X1 U3740 ( .A1(n38501), .A2(n37593), .B1(n38761), .B2(n38498), .ZN(
        n8766) );
  OAI22_X1 U3741 ( .A1(n38501), .A2(n37594), .B1(n38768), .B2(n38498), .ZN(
        n8767) );
  OAI22_X1 U3742 ( .A1(n38501), .A2(n37595), .B1(n38775), .B2(n38498), .ZN(
        n8768) );
  OAI22_X1 U3743 ( .A1(n38501), .A2(n37596), .B1(n38782), .B2(n38498), .ZN(
        n8769) );
  OAI22_X1 U3744 ( .A1(n38502), .A2(n37597), .B1(n38789), .B2(n38498), .ZN(
        n8770) );
  OAI22_X1 U3745 ( .A1(n38502), .A2(n37598), .B1(n38796), .B2(n3236), .ZN(
        n8771) );
  OAI22_X1 U3746 ( .A1(n38502), .A2(n37599), .B1(n38803), .B2(n38498), .ZN(
        n8772) );
  OAI22_X1 U3747 ( .A1(n38502), .A2(n37600), .B1(n38810), .B2(n3236), .ZN(
        n8773) );
  OAI22_X1 U3748 ( .A1(n38502), .A2(n37601), .B1(n38817), .B2(n3236), .ZN(
        n8774) );
  OAI22_X1 U3749 ( .A1(n38503), .A2(n37602), .B1(n38824), .B2(n3236), .ZN(
        n8775) );
  OAI22_X1 U3750 ( .A1(n38503), .A2(n37603), .B1(n38831), .B2(n3236), .ZN(
        n8776) );
  OAI22_X1 U3751 ( .A1(n38503), .A2(n37604), .B1(n38838), .B2(n38498), .ZN(
        n8777) );
  OAI22_X1 U3752 ( .A1(n38503), .A2(n37605), .B1(n38845), .B2(n3236), .ZN(
        n8778) );
  OAI22_X1 U3753 ( .A1(n38503), .A2(n37606), .B1(n38852), .B2(n3236), .ZN(
        n8779) );
  OAI22_X1 U3754 ( .A1(n38504), .A2(n37607), .B1(n38859), .B2(n3236), .ZN(
        n8780) );
  OAI22_X1 U3755 ( .A1(n38504), .A2(n37608), .B1(n38866), .B2(n38498), .ZN(
        n8781) );
  OAI22_X1 U3756 ( .A1(n38504), .A2(n37609), .B1(n38873), .B2(n3236), .ZN(
        n8782) );
  OAI22_X1 U3757 ( .A1(n38504), .A2(n37610), .B1(n38880), .B2(n38498), .ZN(
        n8783) );
  OAI22_X1 U3758 ( .A1(n38504), .A2(n37611), .B1(n38887), .B2(n3236), .ZN(
        n8784) );
  OAI22_X1 U3759 ( .A1(n38505), .A2(n37612), .B1(n38894), .B2(n38498), .ZN(
        n8785) );
  OAI22_X1 U3760 ( .A1(n38505), .A2(n37613), .B1(n38901), .B2(n3236), .ZN(
        n8786) );
  OAI22_X1 U3761 ( .A1(n38547), .A2(n37454), .B1(n38684), .B2(n38546), .ZN(
        n8883) );
  OAI22_X1 U3762 ( .A1(n38547), .A2(n37455), .B1(n38691), .B2(n38546), .ZN(
        n8884) );
  OAI22_X1 U3763 ( .A1(n38547), .A2(n37456), .B1(n38698), .B2(n38546), .ZN(
        n8885) );
  OAI22_X1 U3764 ( .A1(n38547), .A2(n37457), .B1(n38705), .B2(n38546), .ZN(
        n8886) );
  OAI22_X1 U3765 ( .A1(n38547), .A2(n37458), .B1(n38712), .B2(n38546), .ZN(
        n8887) );
  OAI22_X1 U3766 ( .A1(n38548), .A2(n37459), .B1(n38719), .B2(n38546), .ZN(
        n8888) );
  OAI22_X1 U3767 ( .A1(n38548), .A2(n37460), .B1(n38726), .B2(n38546), .ZN(
        n8889) );
  OAI22_X1 U3768 ( .A1(n38548), .A2(n37461), .B1(n38733), .B2(n38546), .ZN(
        n8890) );
  OAI22_X1 U3769 ( .A1(n38548), .A2(n37462), .B1(n38740), .B2(n38546), .ZN(
        n8891) );
  OAI22_X1 U3770 ( .A1(n38548), .A2(n37463), .B1(n38747), .B2(n38546), .ZN(
        n8892) );
  OAI22_X1 U3771 ( .A1(n38549), .A2(n37464), .B1(n38754), .B2(n38546), .ZN(
        n8893) );
  OAI22_X1 U3772 ( .A1(n38549), .A2(n37465), .B1(n38761), .B2(n38546), .ZN(
        n8894) );
  OAI22_X1 U3773 ( .A1(n38549), .A2(n37466), .B1(n38768), .B2(n38546), .ZN(
        n8895) );
  OAI22_X1 U3774 ( .A1(n38549), .A2(n37467), .B1(n38775), .B2(n38546), .ZN(
        n8896) );
  OAI22_X1 U3775 ( .A1(n38549), .A2(n37468), .B1(n38782), .B2(n38546), .ZN(
        n8897) );
  OAI22_X1 U3776 ( .A1(n38550), .A2(n37469), .B1(n38789), .B2(n38546), .ZN(
        n8898) );
  OAI22_X1 U3777 ( .A1(n38550), .A2(n37470), .B1(n38796), .B2(n3096), .ZN(
        n8899) );
  OAI22_X1 U3778 ( .A1(n38550), .A2(n37471), .B1(n38803), .B2(n38546), .ZN(
        n8900) );
  OAI22_X1 U3779 ( .A1(n38550), .A2(n37472), .B1(n38810), .B2(n3096), .ZN(
        n8901) );
  OAI22_X1 U3780 ( .A1(n38550), .A2(n37473), .B1(n38817), .B2(n3096), .ZN(
        n8902) );
  OAI22_X1 U3781 ( .A1(n38551), .A2(n37474), .B1(n38824), .B2(n3096), .ZN(
        n8903) );
  OAI22_X1 U3782 ( .A1(n38551), .A2(n37475), .B1(n38831), .B2(n3096), .ZN(
        n8904) );
  OAI22_X1 U3783 ( .A1(n38551), .A2(n37476), .B1(n38838), .B2(n38546), .ZN(
        n8905) );
  OAI22_X1 U3784 ( .A1(n38551), .A2(n37477), .B1(n38845), .B2(n3096), .ZN(
        n8906) );
  OAI22_X1 U3785 ( .A1(n38551), .A2(n37478), .B1(n38852), .B2(n3096), .ZN(
        n8907) );
  OAI22_X1 U3786 ( .A1(n38552), .A2(n37479), .B1(n38859), .B2(n3096), .ZN(
        n8908) );
  OAI22_X1 U3787 ( .A1(n38552), .A2(n37480), .B1(n38866), .B2(n38546), .ZN(
        n8909) );
  OAI22_X1 U3788 ( .A1(n38552), .A2(n37481), .B1(n38873), .B2(n3096), .ZN(
        n8910) );
  OAI22_X1 U3789 ( .A1(n38552), .A2(n37482), .B1(n38880), .B2(n38546), .ZN(
        n8911) );
  OAI22_X1 U3790 ( .A1(n38552), .A2(n37483), .B1(n38887), .B2(n3096), .ZN(
        n8912) );
  OAI22_X1 U3791 ( .A1(n38553), .A2(n37484), .B1(n38894), .B2(n38546), .ZN(
        n8913) );
  OAI22_X1 U3792 ( .A1(n38553), .A2(n37485), .B1(n38901), .B2(n3096), .ZN(
        n8914) );
  OAI22_X1 U3793 ( .A1(n38559), .A2(n37614), .B1(n38684), .B2(n38558), .ZN(
        n8915) );
  OAI22_X1 U3794 ( .A1(n38559), .A2(n37615), .B1(n38691), .B2(n38558), .ZN(
        n8916) );
  OAI22_X1 U3795 ( .A1(n38559), .A2(n37616), .B1(n38698), .B2(n38558), .ZN(
        n8917) );
  OAI22_X1 U3796 ( .A1(n38559), .A2(n37617), .B1(n38705), .B2(n38558), .ZN(
        n8918) );
  OAI22_X1 U3797 ( .A1(n38559), .A2(n37618), .B1(n38712), .B2(n38558), .ZN(
        n8919) );
  OAI22_X1 U3798 ( .A1(n38560), .A2(n37619), .B1(n38719), .B2(n38558), .ZN(
        n8920) );
  OAI22_X1 U3799 ( .A1(n38560), .A2(n37620), .B1(n38726), .B2(n38558), .ZN(
        n8921) );
  OAI22_X1 U3800 ( .A1(n38560), .A2(n37621), .B1(n38733), .B2(n38558), .ZN(
        n8922) );
  OAI22_X1 U3801 ( .A1(n38560), .A2(n37622), .B1(n38740), .B2(n38558), .ZN(
        n8923) );
  OAI22_X1 U3802 ( .A1(n38560), .A2(n37623), .B1(n38747), .B2(n38558), .ZN(
        n8924) );
  OAI22_X1 U3803 ( .A1(n38561), .A2(n37624), .B1(n38754), .B2(n38558), .ZN(
        n8925) );
  OAI22_X1 U3804 ( .A1(n38561), .A2(n37625), .B1(n38761), .B2(n38558), .ZN(
        n8926) );
  OAI22_X1 U3805 ( .A1(n38561), .A2(n37626), .B1(n38768), .B2(n38558), .ZN(
        n8927) );
  OAI22_X1 U3806 ( .A1(n38561), .A2(n37627), .B1(n38775), .B2(n38558), .ZN(
        n8928) );
  OAI22_X1 U3807 ( .A1(n38561), .A2(n37628), .B1(n38782), .B2(n38558), .ZN(
        n8929) );
  OAI22_X1 U3808 ( .A1(n38562), .A2(n37629), .B1(n38789), .B2(n38558), .ZN(
        n8930) );
  OAI22_X1 U3809 ( .A1(n38562), .A2(n37630), .B1(n38796), .B2(n3061), .ZN(
        n8931) );
  OAI22_X1 U3810 ( .A1(n38562), .A2(n37631), .B1(n38803), .B2(n38558), .ZN(
        n8932) );
  OAI22_X1 U3811 ( .A1(n38562), .A2(n37632), .B1(n38810), .B2(n3061), .ZN(
        n8933) );
  OAI22_X1 U3812 ( .A1(n38562), .A2(n37633), .B1(n38817), .B2(n3061), .ZN(
        n8934) );
  OAI22_X1 U3813 ( .A1(n38563), .A2(n37634), .B1(n38824), .B2(n3061), .ZN(
        n8935) );
  OAI22_X1 U3814 ( .A1(n38563), .A2(n37635), .B1(n38831), .B2(n3061), .ZN(
        n8936) );
  OAI22_X1 U3815 ( .A1(n38563), .A2(n37636), .B1(n38838), .B2(n38558), .ZN(
        n8937) );
  OAI22_X1 U3816 ( .A1(n38563), .A2(n37637), .B1(n38845), .B2(n3061), .ZN(
        n8938) );
  OAI22_X1 U3817 ( .A1(n38563), .A2(n37638), .B1(n38852), .B2(n3061), .ZN(
        n8939) );
  OAI22_X1 U3818 ( .A1(n38564), .A2(n37639), .B1(n38859), .B2(n3061), .ZN(
        n8940) );
  OAI22_X1 U3819 ( .A1(n38564), .A2(n37640), .B1(n38866), .B2(n38558), .ZN(
        n8941) );
  OAI22_X1 U3820 ( .A1(n38564), .A2(n37641), .B1(n38873), .B2(n3061), .ZN(
        n8942) );
  OAI22_X1 U3821 ( .A1(n38564), .A2(n37642), .B1(n38880), .B2(n38558), .ZN(
        n8943) );
  OAI22_X1 U3822 ( .A1(n38564), .A2(n37643), .B1(n38887), .B2(n3061), .ZN(
        n8944) );
  OAI22_X1 U3823 ( .A1(n38565), .A2(n37644), .B1(n38894), .B2(n38558), .ZN(
        n8945) );
  OAI22_X1 U3824 ( .A1(n38565), .A2(n37645), .B1(n38901), .B2(n3061), .ZN(
        n8946) );
  OAI22_X1 U3825 ( .A1(n38607), .A2(n37486), .B1(n38684), .B2(n38606), .ZN(
        n9043) );
  OAI22_X1 U3826 ( .A1(n38607), .A2(n37487), .B1(n38691), .B2(n38606), .ZN(
        n9044) );
  OAI22_X1 U3827 ( .A1(n38607), .A2(n37488), .B1(n38698), .B2(n38606), .ZN(
        n9045) );
  OAI22_X1 U3828 ( .A1(n38607), .A2(n37489), .B1(n38705), .B2(n38606), .ZN(
        n9046) );
  OAI22_X1 U3829 ( .A1(n38607), .A2(n37490), .B1(n38712), .B2(n38606), .ZN(
        n9047) );
  OAI22_X1 U3830 ( .A1(n38608), .A2(n37491), .B1(n38719), .B2(n38606), .ZN(
        n9048) );
  OAI22_X1 U3831 ( .A1(n38608), .A2(n37492), .B1(n38726), .B2(n38606), .ZN(
        n9049) );
  OAI22_X1 U3832 ( .A1(n38608), .A2(n37493), .B1(n38733), .B2(n38606), .ZN(
        n9050) );
  OAI22_X1 U3833 ( .A1(n38608), .A2(n37494), .B1(n38740), .B2(n38606), .ZN(
        n9051) );
  OAI22_X1 U3834 ( .A1(n38608), .A2(n37495), .B1(n38747), .B2(n38606), .ZN(
        n9052) );
  OAI22_X1 U3835 ( .A1(n38609), .A2(n37496), .B1(n38754), .B2(n38606), .ZN(
        n9053) );
  OAI22_X1 U3836 ( .A1(n38609), .A2(n37497), .B1(n38761), .B2(n38606), .ZN(
        n9054) );
  OAI22_X1 U3837 ( .A1(n38609), .A2(n37498), .B1(n38768), .B2(n38606), .ZN(
        n9055) );
  OAI22_X1 U3838 ( .A1(n38609), .A2(n37499), .B1(n38775), .B2(n38606), .ZN(
        n9056) );
  OAI22_X1 U3839 ( .A1(n38609), .A2(n37500), .B1(n38782), .B2(n38606), .ZN(
        n9057) );
  OAI22_X1 U3840 ( .A1(n38610), .A2(n37501), .B1(n38789), .B2(n38606), .ZN(
        n9058) );
  OAI22_X1 U3841 ( .A1(n38610), .A2(n37502), .B1(n38796), .B2(n2921), .ZN(
        n9059) );
  OAI22_X1 U3842 ( .A1(n38610), .A2(n37503), .B1(n38803), .B2(n38606), .ZN(
        n9060) );
  OAI22_X1 U3843 ( .A1(n38610), .A2(n37504), .B1(n38810), .B2(n2921), .ZN(
        n9061) );
  OAI22_X1 U3844 ( .A1(n38610), .A2(n37505), .B1(n38817), .B2(n2921), .ZN(
        n9062) );
  OAI22_X1 U3845 ( .A1(n38611), .A2(n37506), .B1(n38824), .B2(n2921), .ZN(
        n9063) );
  OAI22_X1 U3846 ( .A1(n38611), .A2(n37507), .B1(n38831), .B2(n2921), .ZN(
        n9064) );
  OAI22_X1 U3847 ( .A1(n38611), .A2(n37508), .B1(n38838), .B2(n38606), .ZN(
        n9065) );
  OAI22_X1 U3848 ( .A1(n38611), .A2(n37509), .B1(n38845), .B2(n2921), .ZN(
        n9066) );
  OAI22_X1 U3849 ( .A1(n38611), .A2(n37510), .B1(n38852), .B2(n2921), .ZN(
        n9067) );
  OAI22_X1 U3850 ( .A1(n38612), .A2(n37511), .B1(n38859), .B2(n2921), .ZN(
        n9068) );
  OAI22_X1 U3851 ( .A1(n38612), .A2(n37512), .B1(n38866), .B2(n38606), .ZN(
        n9069) );
  OAI22_X1 U3852 ( .A1(n38612), .A2(n37513), .B1(n38873), .B2(n2921), .ZN(
        n9070) );
  OAI22_X1 U3853 ( .A1(n38612), .A2(n37514), .B1(n38880), .B2(n38606), .ZN(
        n9071) );
  OAI22_X1 U3854 ( .A1(n38612), .A2(n37515), .B1(n38887), .B2(n2921), .ZN(
        n9072) );
  OAI22_X1 U3855 ( .A1(n38613), .A2(n37516), .B1(n38894), .B2(n38606), .ZN(
        n9073) );
  OAI22_X1 U3856 ( .A1(n38613), .A2(n37517), .B1(n38901), .B2(n2921), .ZN(
        n9074) );
  OAI22_X1 U3857 ( .A1(n38619), .A2(n37646), .B1(n38684), .B2(n38618), .ZN(
        n9075) );
  OAI22_X1 U3858 ( .A1(n38619), .A2(n37647), .B1(n38691), .B2(n38618), .ZN(
        n9076) );
  OAI22_X1 U3859 ( .A1(n38619), .A2(n37648), .B1(n38698), .B2(n38618), .ZN(
        n9077) );
  OAI22_X1 U3860 ( .A1(n38619), .A2(n37649), .B1(n38705), .B2(n38618), .ZN(
        n9078) );
  OAI22_X1 U3861 ( .A1(n38619), .A2(n37650), .B1(n38712), .B2(n38618), .ZN(
        n9079) );
  OAI22_X1 U3862 ( .A1(n38620), .A2(n37651), .B1(n38719), .B2(n38618), .ZN(
        n9080) );
  OAI22_X1 U3863 ( .A1(n38620), .A2(n37652), .B1(n38726), .B2(n38618), .ZN(
        n9081) );
  OAI22_X1 U3864 ( .A1(n38620), .A2(n37653), .B1(n38733), .B2(n38618), .ZN(
        n9082) );
  OAI22_X1 U3865 ( .A1(n38620), .A2(n37654), .B1(n38740), .B2(n38618), .ZN(
        n9083) );
  OAI22_X1 U3866 ( .A1(n38620), .A2(n37655), .B1(n38747), .B2(n38618), .ZN(
        n9084) );
  OAI22_X1 U3867 ( .A1(n38621), .A2(n37656), .B1(n38754), .B2(n38618), .ZN(
        n9085) );
  OAI22_X1 U3868 ( .A1(n38621), .A2(n37657), .B1(n38761), .B2(n38618), .ZN(
        n9086) );
  OAI22_X1 U3869 ( .A1(n38621), .A2(n37658), .B1(n38768), .B2(n38618), .ZN(
        n9087) );
  OAI22_X1 U3870 ( .A1(n38621), .A2(n37659), .B1(n38775), .B2(n38618), .ZN(
        n9088) );
  OAI22_X1 U3871 ( .A1(n38621), .A2(n37660), .B1(n38782), .B2(n38618), .ZN(
        n9089) );
  OAI22_X1 U3872 ( .A1(n38622), .A2(n37661), .B1(n38789), .B2(n38618), .ZN(
        n9090) );
  OAI22_X1 U3873 ( .A1(n38622), .A2(n37662), .B1(n38796), .B2(n2886), .ZN(
        n9091) );
  OAI22_X1 U3874 ( .A1(n38622), .A2(n37663), .B1(n38803), .B2(n38618), .ZN(
        n9092) );
  OAI22_X1 U3875 ( .A1(n38622), .A2(n37664), .B1(n38810), .B2(n2886), .ZN(
        n9093) );
  OAI22_X1 U3876 ( .A1(n38622), .A2(n37665), .B1(n38817), .B2(n2886), .ZN(
        n9094) );
  OAI22_X1 U3877 ( .A1(n38623), .A2(n37666), .B1(n38824), .B2(n2886), .ZN(
        n9095) );
  OAI22_X1 U3878 ( .A1(n38623), .A2(n37667), .B1(n38831), .B2(n2886), .ZN(
        n9096) );
  OAI22_X1 U3879 ( .A1(n38623), .A2(n37668), .B1(n38838), .B2(n38618), .ZN(
        n9097) );
  OAI22_X1 U3880 ( .A1(n38623), .A2(n37669), .B1(n38845), .B2(n2886), .ZN(
        n9098) );
  OAI22_X1 U3881 ( .A1(n38623), .A2(n37670), .B1(n38852), .B2(n2886), .ZN(
        n9099) );
  OAI22_X1 U3882 ( .A1(n38624), .A2(n37671), .B1(n38859), .B2(n2886), .ZN(
        n9100) );
  OAI22_X1 U3883 ( .A1(n38624), .A2(n37672), .B1(n38866), .B2(n38618), .ZN(
        n9101) );
  OAI22_X1 U3884 ( .A1(n38624), .A2(n37673), .B1(n38873), .B2(n2886), .ZN(
        n9102) );
  OAI22_X1 U3885 ( .A1(n38624), .A2(n37674), .B1(n38880), .B2(n38618), .ZN(
        n9103) );
  OAI22_X1 U3886 ( .A1(n38624), .A2(n37675), .B1(n38887), .B2(n2886), .ZN(
        n9104) );
  OAI22_X1 U3887 ( .A1(n38625), .A2(n37676), .B1(n38894), .B2(n38618), .ZN(
        n9105) );
  OAI22_X1 U3888 ( .A1(n38625), .A2(n37677), .B1(n38901), .B2(n2886), .ZN(
        n9106) );
  OAI22_X1 U3889 ( .A1(n38667), .A2(n37518), .B1(n38684), .B2(n38666), .ZN(
        n9203) );
  OAI22_X1 U3890 ( .A1(n38667), .A2(n37519), .B1(n38691), .B2(n38666), .ZN(
        n9204) );
  OAI22_X1 U3891 ( .A1(n38667), .A2(n37520), .B1(n38698), .B2(n38666), .ZN(
        n9205) );
  OAI22_X1 U3892 ( .A1(n38667), .A2(n37521), .B1(n38705), .B2(n38666), .ZN(
        n9206) );
  OAI22_X1 U3893 ( .A1(n38667), .A2(n37522), .B1(n38712), .B2(n38666), .ZN(
        n9207) );
  OAI22_X1 U3894 ( .A1(n38668), .A2(n37523), .B1(n38719), .B2(n38666), .ZN(
        n9208) );
  OAI22_X1 U3895 ( .A1(n38668), .A2(n37524), .B1(n38726), .B2(n38666), .ZN(
        n9209) );
  OAI22_X1 U3896 ( .A1(n38668), .A2(n37525), .B1(n38733), .B2(n38666), .ZN(
        n9210) );
  OAI22_X1 U3897 ( .A1(n38668), .A2(n37526), .B1(n38740), .B2(n38666), .ZN(
        n9211) );
  OAI22_X1 U3898 ( .A1(n38668), .A2(n37527), .B1(n38747), .B2(n38666), .ZN(
        n9212) );
  OAI22_X1 U3899 ( .A1(n38669), .A2(n37528), .B1(n38754), .B2(n38666), .ZN(
        n9213) );
  OAI22_X1 U3900 ( .A1(n38669), .A2(n37529), .B1(n38761), .B2(n38666), .ZN(
        n9214) );
  OAI22_X1 U3901 ( .A1(n38669), .A2(n37530), .B1(n38768), .B2(n38666), .ZN(
        n9215) );
  OAI22_X1 U3902 ( .A1(n38669), .A2(n37531), .B1(n38775), .B2(n38666), .ZN(
        n9216) );
  OAI22_X1 U3903 ( .A1(n38669), .A2(n37532), .B1(n38782), .B2(n38666), .ZN(
        n9217) );
  OAI22_X1 U3904 ( .A1(n38670), .A2(n37533), .B1(n38789), .B2(n38666), .ZN(
        n9218) );
  OAI22_X1 U3905 ( .A1(n38670), .A2(n37534), .B1(n38796), .B2(n2744), .ZN(
        n9219) );
  OAI22_X1 U3906 ( .A1(n38670), .A2(n37535), .B1(n38803), .B2(n38666), .ZN(
        n9220) );
  OAI22_X1 U3907 ( .A1(n38670), .A2(n37536), .B1(n38810), .B2(n2744), .ZN(
        n9221) );
  OAI22_X1 U3908 ( .A1(n38670), .A2(n37537), .B1(n38817), .B2(n2744), .ZN(
        n9222) );
  OAI22_X1 U3909 ( .A1(n38671), .A2(n37538), .B1(n38824), .B2(n2744), .ZN(
        n9223) );
  OAI22_X1 U3910 ( .A1(n38671), .A2(n37539), .B1(n38831), .B2(n2744), .ZN(
        n9224) );
  OAI22_X1 U3911 ( .A1(n38671), .A2(n37540), .B1(n38838), .B2(n38666), .ZN(
        n9225) );
  OAI22_X1 U3912 ( .A1(n38671), .A2(n37541), .B1(n38845), .B2(n2744), .ZN(
        n9226) );
  OAI22_X1 U3913 ( .A1(n38671), .A2(n37542), .B1(n38852), .B2(n2744), .ZN(
        n9227) );
  OAI22_X1 U3914 ( .A1(n38672), .A2(n37543), .B1(n38859), .B2(n2744), .ZN(
        n9228) );
  OAI22_X1 U3915 ( .A1(n38672), .A2(n37544), .B1(n38866), .B2(n38666), .ZN(
        n9229) );
  OAI22_X1 U3916 ( .A1(n38672), .A2(n37545), .B1(n38873), .B2(n2744), .ZN(
        n9230) );
  OAI22_X1 U3917 ( .A1(n38672), .A2(n37546), .B1(n38880), .B2(n38666), .ZN(
        n9231) );
  OAI22_X1 U3918 ( .A1(n38672), .A2(n37547), .B1(n38887), .B2(n2744), .ZN(
        n9232) );
  OAI22_X1 U3919 ( .A1(n38673), .A2(n37548), .B1(n38894), .B2(n38666), .ZN(
        n9233) );
  OAI22_X1 U3920 ( .A1(n38673), .A2(n37549), .B1(n38901), .B2(n2744), .ZN(
        n9234) );
  OAI22_X1 U3921 ( .A1(n37804), .A2(n37550), .B1(n37796), .B2(n38684), .ZN(
        n6676) );
  OAI22_X1 U3922 ( .A1(n37804), .A2(n37551), .B1(n37796), .B2(n38691), .ZN(
        n6678) );
  OAI22_X1 U3923 ( .A1(n37803), .A2(n37552), .B1(n37796), .B2(n38698), .ZN(
        n6680) );
  OAI22_X1 U3924 ( .A1(n37803), .A2(n37553), .B1(n37796), .B2(n38705), .ZN(
        n6682) );
  OAI22_X1 U3925 ( .A1(n37803), .A2(n37554), .B1(n37796), .B2(n38712), .ZN(
        n6684) );
  OAI22_X1 U3926 ( .A1(n37803), .A2(n37555), .B1(n37796), .B2(n38719), .ZN(
        n6686) );
  OAI22_X1 U3927 ( .A1(n37803), .A2(n37556), .B1(n37796), .B2(n38726), .ZN(
        n6688) );
  OAI22_X1 U3928 ( .A1(n37802), .A2(n37557), .B1(n37796), .B2(n38733), .ZN(
        n6690) );
  OAI22_X1 U3929 ( .A1(n37802), .A2(n37558), .B1(n37796), .B2(n38740), .ZN(
        n6692) );
  OAI22_X1 U3930 ( .A1(n37802), .A2(n37559), .B1(n37796), .B2(n38747), .ZN(
        n6694) );
  OAI22_X1 U3931 ( .A1(n37802), .A2(n37560), .B1(n37796), .B2(n38754), .ZN(
        n6696) );
  OAI22_X1 U3932 ( .A1(n37802), .A2(n37561), .B1(n37796), .B2(n38761), .ZN(
        n6698) );
  OAI22_X1 U3933 ( .A1(n37801), .A2(n37562), .B1(n37797), .B2(n38768), .ZN(
        n6700) );
  OAI22_X1 U3934 ( .A1(n37801), .A2(n37563), .B1(n37797), .B2(n38775), .ZN(
        n6702) );
  OAI22_X1 U3935 ( .A1(n37801), .A2(n37564), .B1(n37797), .B2(n38782), .ZN(
        n6704) );
  OAI22_X1 U3936 ( .A1(n37801), .A2(n37565), .B1(n37797), .B2(n38789), .ZN(
        n6706) );
  OAI22_X1 U3937 ( .A1(n37801), .A2(n37566), .B1(n37797), .B2(n38796), .ZN(
        n6708) );
  OAI22_X1 U3938 ( .A1(n37800), .A2(n37567), .B1(n37797), .B2(n38803), .ZN(
        n6710) );
  OAI22_X1 U3939 ( .A1(n37800), .A2(n37568), .B1(n37797), .B2(n38810), .ZN(
        n6712) );
  OAI22_X1 U3940 ( .A1(n37800), .A2(n37569), .B1(n37797), .B2(n38817), .ZN(
        n6714) );
  OAI22_X1 U3941 ( .A1(n37800), .A2(n37570), .B1(n37797), .B2(n38824), .ZN(
        n6716) );
  OAI22_X1 U3942 ( .A1(n37800), .A2(n37571), .B1(n37797), .B2(n38831), .ZN(
        n6718) );
  OAI22_X1 U3943 ( .A1(n37799), .A2(n37572), .B1(n37797), .B2(n38838), .ZN(
        n6720) );
  OAI22_X1 U3944 ( .A1(n37799), .A2(n37573), .B1(n37797), .B2(n38845), .ZN(
        n6722) );
  OAI22_X1 U3945 ( .A1(n37799), .A2(n37574), .B1(n37796), .B2(n38852), .ZN(
        n6724) );
  OAI22_X1 U3946 ( .A1(n37799), .A2(n37575), .B1(n37797), .B2(n38859), .ZN(
        n6726) );
  OAI22_X1 U3947 ( .A1(n37799), .A2(n37576), .B1(n37796), .B2(n38866), .ZN(
        n6728) );
  OAI22_X1 U3948 ( .A1(n37798), .A2(n37577), .B1(n37797), .B2(n38873), .ZN(
        n6730) );
  OAI22_X1 U3949 ( .A1(n37798), .A2(n37578), .B1(n37796), .B2(n38880), .ZN(
        n6732) );
  OAI22_X1 U3950 ( .A1(n37798), .A2(n37579), .B1(n37797), .B2(n38887), .ZN(
        n6734) );
  OAI22_X1 U3951 ( .A1(n37798), .A2(n37580), .B1(n37796), .B2(n38894), .ZN(
        n6736) );
  OAI22_X1 U3952 ( .A1(n37798), .A2(n37581), .B1(n37797), .B2(n38901), .ZN(
        n6738) );
  OAI22_X1 U3953 ( .A1(n38903), .A2(n37678), .B1(n38902), .B2(n38684), .ZN(
        n9235) );
  OAI22_X1 U3954 ( .A1(n38903), .A2(n37679), .B1(n38902), .B2(n38691), .ZN(
        n9236) );
  OAI22_X1 U3955 ( .A1(n38903), .A2(n37680), .B1(n38902), .B2(n38698), .ZN(
        n9237) );
  OAI22_X1 U3956 ( .A1(n38903), .A2(n37681), .B1(n38902), .B2(n38705), .ZN(
        n9238) );
  OAI22_X1 U3957 ( .A1(n38903), .A2(n37682), .B1(n38902), .B2(n38712), .ZN(
        n9239) );
  OAI22_X1 U3958 ( .A1(n38904), .A2(n37683), .B1(n38902), .B2(n38719), .ZN(
        n9240) );
  OAI22_X1 U3959 ( .A1(n38904), .A2(n37684), .B1(n38902), .B2(n38726), .ZN(
        n9241) );
  OAI22_X1 U3960 ( .A1(n38904), .A2(n37685), .B1(n38902), .B2(n38733), .ZN(
        n9242) );
  OAI22_X1 U3961 ( .A1(n38904), .A2(n37686), .B1(n38902), .B2(n38740), .ZN(
        n9243) );
  OAI22_X1 U3962 ( .A1(n38904), .A2(n37687), .B1(n38902), .B2(n38747), .ZN(
        n9244) );
  OAI22_X1 U3963 ( .A1(n38905), .A2(n37688), .B1(n38902), .B2(n38754), .ZN(
        n9245) );
  OAI22_X1 U3964 ( .A1(n38905), .A2(n37689), .B1(n38902), .B2(n38761), .ZN(
        n9246) );
  OAI22_X1 U3965 ( .A1(n38905), .A2(n37690), .B1(n38902), .B2(n38768), .ZN(
        n9247) );
  OAI22_X1 U3966 ( .A1(n38905), .A2(n37691), .B1(n2676), .B2(n38775), .ZN(
        n9248) );
  OAI22_X1 U3967 ( .A1(n38905), .A2(n37692), .B1(n2676), .B2(n38782), .ZN(
        n9249) );
  OAI22_X1 U3968 ( .A1(n38906), .A2(n37693), .B1(n2676), .B2(n38789), .ZN(
        n9250) );
  OAI22_X1 U3969 ( .A1(n38906), .A2(n37694), .B1(n2676), .B2(n38796), .ZN(
        n9251) );
  OAI22_X1 U3970 ( .A1(n38906), .A2(n37695), .B1(n2676), .B2(n38803), .ZN(
        n9252) );
  OAI22_X1 U3971 ( .A1(n38906), .A2(n37696), .B1(n2676), .B2(n38810), .ZN(
        n9253) );
  OAI22_X1 U3972 ( .A1(n38906), .A2(n37697), .B1(n2676), .B2(n38817), .ZN(
        n9254) );
  OAI22_X1 U3973 ( .A1(n38907), .A2(n37698), .B1(n2676), .B2(n38824), .ZN(
        n9255) );
  OAI22_X1 U3974 ( .A1(n38907), .A2(n37699), .B1(n2676), .B2(n38831), .ZN(
        n9256) );
  OAI22_X1 U3975 ( .A1(n38907), .A2(n37700), .B1(n38902), .B2(n38838), .ZN(
        n9257) );
  OAI22_X1 U3976 ( .A1(n38907), .A2(n37701), .B1(n38902), .B2(n38845), .ZN(
        n9258) );
  OAI22_X1 U3977 ( .A1(n38907), .A2(n37702), .B1(n2676), .B2(n38852), .ZN(
        n9259) );
  OAI22_X1 U3978 ( .A1(n38908), .A2(n37703), .B1(n38902), .B2(n38859), .ZN(
        n9260) );
  OAI22_X1 U3979 ( .A1(n38908), .A2(n37704), .B1(n38902), .B2(n38866), .ZN(
        n9261) );
  OAI22_X1 U3980 ( .A1(n38908), .A2(n37705), .B1(n38902), .B2(n38873), .ZN(
        n9262) );
  OAI22_X1 U3981 ( .A1(n38908), .A2(n37706), .B1(n38902), .B2(n38880), .ZN(
        n9263) );
  OAI22_X1 U3982 ( .A1(n38908), .A2(n37707), .B1(n38902), .B2(n38887), .ZN(
        n9264) );
  OAI22_X1 U3983 ( .A1(n38909), .A2(n37708), .B1(n38902), .B2(n38894), .ZN(
        n9265) );
  OAI22_X1 U3984 ( .A1(n38909), .A2(n37709), .B1(n2676), .B2(n38901), .ZN(
        n9266) );
  INV_X1 U3985 ( .A(ENABLE), .ZN(n9631) );
  OAI22_X1 U3986 ( .A1(n37810), .A2(n38851), .B1(n5474), .B2(n37070), .ZN(
        n6763) );
  OAI22_X1 U3987 ( .A1(n37811), .A2(n38858), .B1(n5474), .B2(n37071), .ZN(
        n6764) );
  OAI22_X1 U3988 ( .A1(n37811), .A2(n38865), .B1(n5474), .B2(n37072), .ZN(
        n6765) );
  OAI22_X1 U3989 ( .A1(n37811), .A2(n38872), .B1(n37805), .B2(n37073), .ZN(
        n6766) );
  OAI22_X1 U3990 ( .A1(n37811), .A2(n38879), .B1(n37805), .B2(n37074), .ZN(
        n6767) );
  OAI22_X1 U3991 ( .A1(n37811), .A2(n38886), .B1(n37805), .B2(n37075), .ZN(
        n6768) );
  OAI22_X1 U3992 ( .A1(n37812), .A2(n38893), .B1(n37805), .B2(n37076), .ZN(
        n6769) );
  OAI22_X1 U3993 ( .A1(n37812), .A2(n38900), .B1(n5474), .B2(n37077), .ZN(
        n6770) );
  OAI22_X1 U3994 ( .A1(n37855), .A2(n38851), .B1(n5334), .B2(n36686), .ZN(
        n6891) );
  OAI22_X1 U3995 ( .A1(n37856), .A2(n38858), .B1(n5334), .B2(n36687), .ZN(
        n6892) );
  OAI22_X1 U3996 ( .A1(n37856), .A2(n38865), .B1(n5334), .B2(n36688), .ZN(
        n6893) );
  OAI22_X1 U3997 ( .A1(n37856), .A2(n38872), .B1(n37850), .B2(n36689), .ZN(
        n6894) );
  OAI22_X1 U3998 ( .A1(n37856), .A2(n38879), .B1(n37850), .B2(n36690), .ZN(
        n6895) );
  OAI22_X1 U3999 ( .A1(n37856), .A2(n38886), .B1(n37850), .B2(n36691), .ZN(
        n6896) );
  OAI22_X1 U4000 ( .A1(n37857), .A2(n38893), .B1(n37850), .B2(n36692), .ZN(
        n6897) );
  OAI22_X1 U4001 ( .A1(n37857), .A2(n38900), .B1(n5334), .B2(n36693), .ZN(
        n6898) );
  OAI22_X1 U4002 ( .A1(n37864), .A2(n38851), .B1(n5299), .B2(n37078), .ZN(
        n6923) );
  OAI22_X1 U4003 ( .A1(n37865), .A2(n38858), .B1(n5299), .B2(n37079), .ZN(
        n6924) );
  OAI22_X1 U4004 ( .A1(n37865), .A2(n38865), .B1(n5299), .B2(n37080), .ZN(
        n6925) );
  OAI22_X1 U4005 ( .A1(n37865), .A2(n38872), .B1(n37859), .B2(n37081), .ZN(
        n6926) );
  OAI22_X1 U4006 ( .A1(n37865), .A2(n38879), .B1(n37859), .B2(n37082), .ZN(
        n6927) );
  OAI22_X1 U4007 ( .A1(n37865), .A2(n38886), .B1(n37859), .B2(n37083), .ZN(
        n6928) );
  OAI22_X1 U4008 ( .A1(n37866), .A2(n38893), .B1(n37859), .B2(n37084), .ZN(
        n6929) );
  OAI22_X1 U4009 ( .A1(n37866), .A2(n38900), .B1(n5299), .B2(n37085), .ZN(
        n6930) );
  OAI22_X1 U4010 ( .A1(n37909), .A2(n38851), .B1(n5159), .B2(n36694), .ZN(
        n7051) );
  OAI22_X1 U4011 ( .A1(n37910), .A2(n38858), .B1(n5159), .B2(n36695), .ZN(
        n7052) );
  OAI22_X1 U4012 ( .A1(n37910), .A2(n38865), .B1(n5159), .B2(n36696), .ZN(
        n7053) );
  OAI22_X1 U4013 ( .A1(n37910), .A2(n38872), .B1(n37904), .B2(n36697), .ZN(
        n7054) );
  OAI22_X1 U4014 ( .A1(n37910), .A2(n38879), .B1(n37904), .B2(n36698), .ZN(
        n7055) );
  OAI22_X1 U4015 ( .A1(n37910), .A2(n38886), .B1(n37904), .B2(n36699), .ZN(
        n7056) );
  OAI22_X1 U4016 ( .A1(n37911), .A2(n38893), .B1(n37904), .B2(n36700), .ZN(
        n7057) );
  OAI22_X1 U4017 ( .A1(n37911), .A2(n38900), .B1(n5159), .B2(n36701), .ZN(
        n7058) );
  OAI22_X1 U4018 ( .A1(n37918), .A2(n38851), .B1(n5124), .B2(n37086), .ZN(
        n7083) );
  OAI22_X1 U4019 ( .A1(n37919), .A2(n38858), .B1(n5124), .B2(n37087), .ZN(
        n7084) );
  OAI22_X1 U4020 ( .A1(n37919), .A2(n38865), .B1(n5124), .B2(n37088), .ZN(
        n7085) );
  OAI22_X1 U4021 ( .A1(n37919), .A2(n38872), .B1(n37913), .B2(n37089), .ZN(
        n7086) );
  OAI22_X1 U4022 ( .A1(n37919), .A2(n38879), .B1(n37913), .B2(n37090), .ZN(
        n7087) );
  OAI22_X1 U4023 ( .A1(n37919), .A2(n38886), .B1(n37913), .B2(n37091), .ZN(
        n7088) );
  OAI22_X1 U4024 ( .A1(n37920), .A2(n38893), .B1(n37913), .B2(n37092), .ZN(
        n7089) );
  OAI22_X1 U4025 ( .A1(n37920), .A2(n38900), .B1(n5124), .B2(n37093), .ZN(
        n7090) );
  OAI22_X1 U4026 ( .A1(n37963), .A2(n38850), .B1(n4983), .B2(n36702), .ZN(
        n7211) );
  OAI22_X1 U4027 ( .A1(n37964), .A2(n38857), .B1(n4983), .B2(n36703), .ZN(
        n7212) );
  OAI22_X1 U4028 ( .A1(n37964), .A2(n38864), .B1(n4983), .B2(n36704), .ZN(
        n7213) );
  OAI22_X1 U4029 ( .A1(n37964), .A2(n38871), .B1(n37958), .B2(n36705), .ZN(
        n7214) );
  OAI22_X1 U4030 ( .A1(n37964), .A2(n38878), .B1(n37958), .B2(n36706), .ZN(
        n7215) );
  OAI22_X1 U4031 ( .A1(n37964), .A2(n38885), .B1(n37958), .B2(n36707), .ZN(
        n7216) );
  OAI22_X1 U4032 ( .A1(n37965), .A2(n38892), .B1(n37958), .B2(n36708), .ZN(
        n7217) );
  OAI22_X1 U4033 ( .A1(n37965), .A2(n38899), .B1(n4983), .B2(n36709), .ZN(
        n7218) );
  OAI22_X1 U4034 ( .A1(n37996), .A2(n38850), .B1(n4878), .B2(n36710), .ZN(
        n7307) );
  OAI22_X1 U4035 ( .A1(n37997), .A2(n38857), .B1(n4878), .B2(n36711), .ZN(
        n7308) );
  OAI22_X1 U4036 ( .A1(n37997), .A2(n38864), .B1(n4878), .B2(n36712), .ZN(
        n7309) );
  OAI22_X1 U4037 ( .A1(n37997), .A2(n38871), .B1(n37991), .B2(n36713), .ZN(
        n7310) );
  OAI22_X1 U4038 ( .A1(n37997), .A2(n38878), .B1(n37991), .B2(n36714), .ZN(
        n7311) );
  OAI22_X1 U4039 ( .A1(n37997), .A2(n38885), .B1(n37991), .B2(n36715), .ZN(
        n7312) );
  OAI22_X1 U4040 ( .A1(n37998), .A2(n38892), .B1(n37991), .B2(n36716), .ZN(
        n7313) );
  OAI22_X1 U4041 ( .A1(n37998), .A2(n38899), .B1(n4878), .B2(n36717), .ZN(
        n7314) );
  OAI22_X1 U4042 ( .A1(n38017), .A2(n38849), .B1(n4808), .B2(n37094), .ZN(
        n7371) );
  OAI22_X1 U4043 ( .A1(n38018), .A2(n38856), .B1(n4808), .B2(n37095), .ZN(
        n7372) );
  OAI22_X1 U4044 ( .A1(n38018), .A2(n38863), .B1(n4808), .B2(n37096), .ZN(
        n7373) );
  OAI22_X1 U4045 ( .A1(n38018), .A2(n38870), .B1(n38012), .B2(n37097), .ZN(
        n7374) );
  OAI22_X1 U4046 ( .A1(n38018), .A2(n38877), .B1(n38012), .B2(n37098), .ZN(
        n7375) );
  OAI22_X1 U4047 ( .A1(n38018), .A2(n38884), .B1(n38012), .B2(n37099), .ZN(
        n7376) );
  OAI22_X1 U4048 ( .A1(n38019), .A2(n38891), .B1(n38012), .B2(n37100), .ZN(
        n7377) );
  OAI22_X1 U4049 ( .A1(n38019), .A2(n38898), .B1(n4808), .B2(n37101), .ZN(
        n7378) );
  OAI22_X1 U4050 ( .A1(n38050), .A2(n38850), .B1(n4703), .B2(n36718), .ZN(
        n7467) );
  OAI22_X1 U4051 ( .A1(n38051), .A2(n38857), .B1(n4703), .B2(n36719), .ZN(
        n7468) );
  OAI22_X1 U4052 ( .A1(n38051), .A2(n38864), .B1(n4703), .B2(n36720), .ZN(
        n7469) );
  OAI22_X1 U4053 ( .A1(n38051), .A2(n38871), .B1(n38045), .B2(n36721), .ZN(
        n7470) );
  OAI22_X1 U4054 ( .A1(n38051), .A2(n38878), .B1(n38045), .B2(n36722), .ZN(
        n7471) );
  OAI22_X1 U4055 ( .A1(n38051), .A2(n38885), .B1(n38045), .B2(n36723), .ZN(
        n7472) );
  OAI22_X1 U4056 ( .A1(n38052), .A2(n38892), .B1(n38045), .B2(n36724), .ZN(
        n7473) );
  OAI22_X1 U4057 ( .A1(n38052), .A2(n38899), .B1(n4703), .B2(n36725), .ZN(
        n7474) );
  OAI22_X1 U4058 ( .A1(n38071), .A2(n38850), .B1(n4633), .B2(n37102), .ZN(
        n7531) );
  OAI22_X1 U4059 ( .A1(n38072), .A2(n38857), .B1(n4633), .B2(n37103), .ZN(
        n7532) );
  OAI22_X1 U4060 ( .A1(n38072), .A2(n38864), .B1(n4633), .B2(n37104), .ZN(
        n7533) );
  OAI22_X1 U4061 ( .A1(n38072), .A2(n38871), .B1(n38066), .B2(n37105), .ZN(
        n7534) );
  OAI22_X1 U4062 ( .A1(n38072), .A2(n38878), .B1(n38066), .B2(n37106), .ZN(
        n7535) );
  OAI22_X1 U4063 ( .A1(n38072), .A2(n38885), .B1(n38066), .B2(n37107), .ZN(
        n7536) );
  OAI22_X1 U4064 ( .A1(n38073), .A2(n38892), .B1(n38066), .B2(n37108), .ZN(
        n7537) );
  OAI22_X1 U4065 ( .A1(n38073), .A2(n38899), .B1(n4633), .B2(n37109), .ZN(
        n7538) );
  OAI22_X1 U4066 ( .A1(n38104), .A2(n38849), .B1(n4528), .B2(n36726), .ZN(
        n7627) );
  OAI22_X1 U4067 ( .A1(n38105), .A2(n38856), .B1(n4528), .B2(n36727), .ZN(
        n7628) );
  OAI22_X1 U4068 ( .A1(n38105), .A2(n38863), .B1(n4528), .B2(n36728), .ZN(
        n7629) );
  OAI22_X1 U4069 ( .A1(n38105), .A2(n38870), .B1(n38099), .B2(n36729), .ZN(
        n7630) );
  OAI22_X1 U4070 ( .A1(n38105), .A2(n38877), .B1(n38099), .B2(n36730), .ZN(
        n7631) );
  OAI22_X1 U4071 ( .A1(n38105), .A2(n38884), .B1(n38099), .B2(n36731), .ZN(
        n7632) );
  OAI22_X1 U4072 ( .A1(n38106), .A2(n38891), .B1(n38099), .B2(n36732), .ZN(
        n7633) );
  OAI22_X1 U4073 ( .A1(n38106), .A2(n38898), .B1(n4528), .B2(n36733), .ZN(
        n7634) );
  OAI22_X1 U4074 ( .A1(n38125), .A2(n38849), .B1(n4458), .B2(n37110), .ZN(
        n7691) );
  OAI22_X1 U4075 ( .A1(n38126), .A2(n38856), .B1(n4458), .B2(n37111), .ZN(
        n7692) );
  OAI22_X1 U4076 ( .A1(n38126), .A2(n38863), .B1(n4458), .B2(n37112), .ZN(
        n7693) );
  OAI22_X1 U4077 ( .A1(n38126), .A2(n38870), .B1(n38120), .B2(n37113), .ZN(
        n7694) );
  OAI22_X1 U4078 ( .A1(n38126), .A2(n38877), .B1(n38120), .B2(n37114), .ZN(
        n7695) );
  OAI22_X1 U4079 ( .A1(n38126), .A2(n38884), .B1(n38120), .B2(n37115), .ZN(
        n7696) );
  OAI22_X1 U4080 ( .A1(n38127), .A2(n38891), .B1(n38120), .B2(n37116), .ZN(
        n7697) );
  OAI22_X1 U4081 ( .A1(n38127), .A2(n38898), .B1(n4458), .B2(n37117), .ZN(
        n7698) );
  OAI22_X1 U4082 ( .A1(n38158), .A2(n38849), .B1(n4353), .B2(n37118), .ZN(
        n7787) );
  OAI22_X1 U4083 ( .A1(n38159), .A2(n38856), .B1(n4353), .B2(n37119), .ZN(
        n7788) );
  OAI22_X1 U4084 ( .A1(n38159), .A2(n38863), .B1(n4353), .B2(n37120), .ZN(
        n7789) );
  OAI22_X1 U4085 ( .A1(n38159), .A2(n38870), .B1(n38153), .B2(n37121), .ZN(
        n7790) );
  OAI22_X1 U4086 ( .A1(n38159), .A2(n38877), .B1(n38153), .B2(n37122), .ZN(
        n7791) );
  OAI22_X1 U4087 ( .A1(n38159), .A2(n38884), .B1(n38153), .B2(n37123), .ZN(
        n7792) );
  OAI22_X1 U4088 ( .A1(n38160), .A2(n38891), .B1(n38153), .B2(n37124), .ZN(
        n7793) );
  OAI22_X1 U4089 ( .A1(n38160), .A2(n38898), .B1(n4353), .B2(n37125), .ZN(
        n7794) );
  OAI22_X1 U4090 ( .A1(n38191), .A2(n38849), .B1(n4248), .B2(n36734), .ZN(
        n7883) );
  OAI22_X1 U4091 ( .A1(n38192), .A2(n38856), .B1(n4248), .B2(n36735), .ZN(
        n7884) );
  OAI22_X1 U4092 ( .A1(n38192), .A2(n38863), .B1(n4248), .B2(n36736), .ZN(
        n7885) );
  OAI22_X1 U4093 ( .A1(n38192), .A2(n38870), .B1(n38186), .B2(n36737), .ZN(
        n7886) );
  OAI22_X1 U4094 ( .A1(n38192), .A2(n38877), .B1(n38186), .B2(n36738), .ZN(
        n7887) );
  OAI22_X1 U4095 ( .A1(n38192), .A2(n38884), .B1(n38186), .B2(n36739), .ZN(
        n7888) );
  OAI22_X1 U4096 ( .A1(n38193), .A2(n38891), .B1(n38186), .B2(n36740), .ZN(
        n7889) );
  OAI22_X1 U4097 ( .A1(n38193), .A2(n38898), .B1(n4248), .B2(n36741), .ZN(
        n7890) );
  OAI22_X1 U4098 ( .A1(n38212), .A2(n38848), .B1(n4178), .B2(n37126), .ZN(
        n7947) );
  OAI22_X1 U4099 ( .A1(n38213), .A2(n38855), .B1(n4178), .B2(n37127), .ZN(
        n7948) );
  OAI22_X1 U4100 ( .A1(n38213), .A2(n38862), .B1(n4178), .B2(n37128), .ZN(
        n7949) );
  OAI22_X1 U4101 ( .A1(n38213), .A2(n38869), .B1(n38207), .B2(n37129), .ZN(
        n7950) );
  OAI22_X1 U4102 ( .A1(n38213), .A2(n38876), .B1(n38207), .B2(n37130), .ZN(
        n7951) );
  OAI22_X1 U4103 ( .A1(n38213), .A2(n38883), .B1(n38207), .B2(n37131), .ZN(
        n7952) );
  OAI22_X1 U4104 ( .A1(n38214), .A2(n38890), .B1(n38207), .B2(n37132), .ZN(
        n7953) );
  OAI22_X1 U4105 ( .A1(n38214), .A2(n38897), .B1(n4178), .B2(n37133), .ZN(
        n7954) );
  OAI22_X1 U4106 ( .A1(n38245), .A2(n38848), .B1(n4041), .B2(n36742), .ZN(
        n8043) );
  OAI22_X1 U4107 ( .A1(n38246), .A2(n38855), .B1(n4041), .B2(n36743), .ZN(
        n8044) );
  OAI22_X1 U4108 ( .A1(n38246), .A2(n38862), .B1(n4041), .B2(n36744), .ZN(
        n8045) );
  OAI22_X1 U4109 ( .A1(n38246), .A2(n38869), .B1(n38240), .B2(n36745), .ZN(
        n8046) );
  OAI22_X1 U4110 ( .A1(n38246), .A2(n38876), .B1(n38240), .B2(n36746), .ZN(
        n8047) );
  OAI22_X1 U4111 ( .A1(n38246), .A2(n38883), .B1(n38240), .B2(n36747), .ZN(
        n8048) );
  OAI22_X1 U4112 ( .A1(n38247), .A2(n38890), .B1(n38240), .B2(n36748), .ZN(
        n8049) );
  OAI22_X1 U4113 ( .A1(n38247), .A2(n38897), .B1(n4041), .B2(n36749), .ZN(
        n8050) );
  OAI22_X1 U4114 ( .A1(n38266), .A2(n38848), .B1(n3971), .B2(n37134), .ZN(
        n8107) );
  OAI22_X1 U4115 ( .A1(n38267), .A2(n38855), .B1(n3971), .B2(n37135), .ZN(
        n8108) );
  OAI22_X1 U4116 ( .A1(n38267), .A2(n38862), .B1(n3971), .B2(n37136), .ZN(
        n8109) );
  OAI22_X1 U4117 ( .A1(n38267), .A2(n38869), .B1(n38261), .B2(n37137), .ZN(
        n8110) );
  OAI22_X1 U4118 ( .A1(n38267), .A2(n38876), .B1(n38261), .B2(n37138), .ZN(
        n8111) );
  OAI22_X1 U4119 ( .A1(n38267), .A2(n38883), .B1(n38261), .B2(n37139), .ZN(
        n8112) );
  OAI22_X1 U4120 ( .A1(n38268), .A2(n38890), .B1(n38261), .B2(n37140), .ZN(
        n8113) );
  OAI22_X1 U4121 ( .A1(n38268), .A2(n38897), .B1(n3971), .B2(n37141), .ZN(
        n8114) );
  OAI22_X1 U4122 ( .A1(n38299), .A2(n38848), .B1(n3866), .B2(n36750), .ZN(
        n8203) );
  OAI22_X1 U4123 ( .A1(n38300), .A2(n38855), .B1(n3866), .B2(n36751), .ZN(
        n8204) );
  OAI22_X1 U4124 ( .A1(n38300), .A2(n38862), .B1(n3866), .B2(n36752), .ZN(
        n8205) );
  OAI22_X1 U4125 ( .A1(n38300), .A2(n38869), .B1(n38294), .B2(n36753), .ZN(
        n8206) );
  OAI22_X1 U4126 ( .A1(n38300), .A2(n38876), .B1(n38294), .B2(n36754), .ZN(
        n8207) );
  OAI22_X1 U4127 ( .A1(n38300), .A2(n38883), .B1(n38294), .B2(n36755), .ZN(
        n8208) );
  OAI22_X1 U4128 ( .A1(n38301), .A2(n38890), .B1(n38294), .B2(n36756), .ZN(
        n8209) );
  OAI22_X1 U4129 ( .A1(n38301), .A2(n38897), .B1(n3866), .B2(n36757), .ZN(
        n8210) );
  OAI22_X1 U4130 ( .A1(n38332), .A2(n38847), .B1(n3761), .B2(n36758), .ZN(
        n8299) );
  OAI22_X1 U4131 ( .A1(n38333), .A2(n38854), .B1(n3761), .B2(n36759), .ZN(
        n8300) );
  OAI22_X1 U4132 ( .A1(n38333), .A2(n38861), .B1(n3761), .B2(n36760), .ZN(
        n8301) );
  OAI22_X1 U4133 ( .A1(n38333), .A2(n38868), .B1(n38327), .B2(n36761), .ZN(
        n8302) );
  OAI22_X1 U4134 ( .A1(n38333), .A2(n38875), .B1(n38327), .B2(n36762), .ZN(
        n8303) );
  OAI22_X1 U4135 ( .A1(n38333), .A2(n38882), .B1(n38327), .B2(n36763), .ZN(
        n8304) );
  OAI22_X1 U4136 ( .A1(n38334), .A2(n38889), .B1(n38327), .B2(n36764), .ZN(
        n8305) );
  OAI22_X1 U4137 ( .A1(n38334), .A2(n38896), .B1(n3761), .B2(n36765), .ZN(
        n8306) );
  OAI22_X1 U4138 ( .A1(n38353), .A2(n38847), .B1(n3691), .B2(n37142), .ZN(
        n8363) );
  OAI22_X1 U4139 ( .A1(n38354), .A2(n38854), .B1(n3691), .B2(n37143), .ZN(
        n8364) );
  OAI22_X1 U4140 ( .A1(n38354), .A2(n38861), .B1(n3691), .B2(n37144), .ZN(
        n8365) );
  OAI22_X1 U4141 ( .A1(n38354), .A2(n38868), .B1(n38348), .B2(n37145), .ZN(
        n8366) );
  OAI22_X1 U4142 ( .A1(n38354), .A2(n38875), .B1(n38348), .B2(n37146), .ZN(
        n8367) );
  OAI22_X1 U4143 ( .A1(n38354), .A2(n38882), .B1(n38348), .B2(n37147), .ZN(
        n8368) );
  OAI22_X1 U4144 ( .A1(n38355), .A2(n38889), .B1(n38348), .B2(n37148), .ZN(
        n8369) );
  OAI22_X1 U4145 ( .A1(n38355), .A2(n38896), .B1(n3691), .B2(n37149), .ZN(
        n8370) );
  OAI22_X1 U4146 ( .A1(n38386), .A2(n38847), .B1(n3586), .B2(n36766), .ZN(
        n8459) );
  OAI22_X1 U4147 ( .A1(n38387), .A2(n38854), .B1(n3586), .B2(n36767), .ZN(
        n8460) );
  OAI22_X1 U4148 ( .A1(n38387), .A2(n38861), .B1(n3586), .B2(n36768), .ZN(
        n8461) );
  OAI22_X1 U4149 ( .A1(n38387), .A2(n38868), .B1(n38381), .B2(n36769), .ZN(
        n8462) );
  OAI22_X1 U4150 ( .A1(n38387), .A2(n38875), .B1(n38381), .B2(n36770), .ZN(
        n8463) );
  OAI22_X1 U4151 ( .A1(n38387), .A2(n38882), .B1(n38381), .B2(n36771), .ZN(
        n8464) );
  OAI22_X1 U4152 ( .A1(n38388), .A2(n38889), .B1(n38381), .B2(n36772), .ZN(
        n8465) );
  OAI22_X1 U4153 ( .A1(n38388), .A2(n38896), .B1(n3586), .B2(n36773), .ZN(
        n8466) );
  OAI22_X1 U4154 ( .A1(n38407), .A2(n38847), .B1(n3516), .B2(n37150), .ZN(
        n8523) );
  OAI22_X1 U4155 ( .A1(n38408), .A2(n38854), .B1(n3516), .B2(n37151), .ZN(
        n8524) );
  OAI22_X1 U4156 ( .A1(n38408), .A2(n38861), .B1(n3516), .B2(n37152), .ZN(
        n8525) );
  OAI22_X1 U4157 ( .A1(n38408), .A2(n38868), .B1(n38402), .B2(n37153), .ZN(
        n8526) );
  OAI22_X1 U4158 ( .A1(n38408), .A2(n38875), .B1(n38402), .B2(n37154), .ZN(
        n8527) );
  OAI22_X1 U4159 ( .A1(n38408), .A2(n38882), .B1(n38402), .B2(n37155), .ZN(
        n8528) );
  OAI22_X1 U4160 ( .A1(n38409), .A2(n38889), .B1(n38402), .B2(n37156), .ZN(
        n8529) );
  OAI22_X1 U4161 ( .A1(n38409), .A2(n38896), .B1(n3516), .B2(n37157), .ZN(
        n8530) );
  OAI22_X1 U4162 ( .A1(n38440), .A2(n38847), .B1(n3411), .B2(n36774), .ZN(
        n8619) );
  OAI22_X1 U4163 ( .A1(n38441), .A2(n38854), .B1(n3411), .B2(n36775), .ZN(
        n8620) );
  OAI22_X1 U4164 ( .A1(n38441), .A2(n38861), .B1(n3411), .B2(n36776), .ZN(
        n8621) );
  OAI22_X1 U4165 ( .A1(n38441), .A2(n38868), .B1(n38435), .B2(n36777), .ZN(
        n8622) );
  OAI22_X1 U4166 ( .A1(n38441), .A2(n38875), .B1(n38435), .B2(n36778), .ZN(
        n8623) );
  OAI22_X1 U4167 ( .A1(n38441), .A2(n38882), .B1(n38435), .B2(n36779), .ZN(
        n8624) );
  OAI22_X1 U4168 ( .A1(n38442), .A2(n38889), .B1(n38435), .B2(n36780), .ZN(
        n8625) );
  OAI22_X1 U4169 ( .A1(n38442), .A2(n38896), .B1(n3411), .B2(n36781), .ZN(
        n8626) );
  OAI22_X1 U4170 ( .A1(n38461), .A2(n38846), .B1(n3341), .B2(n37158), .ZN(
        n8683) );
  OAI22_X1 U4171 ( .A1(n38462), .A2(n38853), .B1(n3341), .B2(n37159), .ZN(
        n8684) );
  OAI22_X1 U4172 ( .A1(n38462), .A2(n38860), .B1(n3341), .B2(n37160), .ZN(
        n8685) );
  OAI22_X1 U4173 ( .A1(n38462), .A2(n38867), .B1(n38456), .B2(n37161), .ZN(
        n8686) );
  OAI22_X1 U4174 ( .A1(n38462), .A2(n38874), .B1(n38456), .B2(n37162), .ZN(
        n8687) );
  OAI22_X1 U4175 ( .A1(n38462), .A2(n38881), .B1(n38456), .B2(n37163), .ZN(
        n8688) );
  OAI22_X1 U4176 ( .A1(n38463), .A2(n38888), .B1(n38456), .B2(n37164), .ZN(
        n8689) );
  OAI22_X1 U4177 ( .A1(n38463), .A2(n38895), .B1(n3341), .B2(n37165), .ZN(
        n8690) );
  OAI22_X1 U4178 ( .A1(n37806), .A2(n38683), .B1(n37805), .B2(n37166), .ZN(
        n6739) );
  OAI22_X1 U4179 ( .A1(n37806), .A2(n38690), .B1(n37805), .B2(n37167), .ZN(
        n6740) );
  OAI22_X1 U4180 ( .A1(n37806), .A2(n38697), .B1(n37805), .B2(n37168), .ZN(
        n6741) );
  OAI22_X1 U4181 ( .A1(n37806), .A2(n38704), .B1(n37805), .B2(n37169), .ZN(
        n6742) );
  OAI22_X1 U4182 ( .A1(n37806), .A2(n38711), .B1(n37805), .B2(n37170), .ZN(
        n6743) );
  OAI22_X1 U4183 ( .A1(n37807), .A2(n38718), .B1(n37805), .B2(n37171), .ZN(
        n6744) );
  OAI22_X1 U4184 ( .A1(n37807), .A2(n38725), .B1(n37805), .B2(n37172), .ZN(
        n6745) );
  OAI22_X1 U4185 ( .A1(n37807), .A2(n38732), .B1(n37805), .B2(n37173), .ZN(
        n6746) );
  OAI22_X1 U4186 ( .A1(n37807), .A2(n38739), .B1(n37805), .B2(n37174), .ZN(
        n6747) );
  OAI22_X1 U4187 ( .A1(n37807), .A2(n38746), .B1(n37805), .B2(n37175), .ZN(
        n6748) );
  OAI22_X1 U4188 ( .A1(n37808), .A2(n38753), .B1(n37805), .B2(n37176), .ZN(
        n6749) );
  OAI22_X1 U4189 ( .A1(n37808), .A2(n38760), .B1(n37805), .B2(n37177), .ZN(
        n6750) );
  OAI22_X1 U4190 ( .A1(n37808), .A2(n38767), .B1(n37805), .B2(n37178), .ZN(
        n6751) );
  OAI22_X1 U4191 ( .A1(n37808), .A2(n38774), .B1(n37805), .B2(n37179), .ZN(
        n6752) );
  OAI22_X1 U4192 ( .A1(n37808), .A2(n38781), .B1(n5474), .B2(n37180), .ZN(
        n6753) );
  OAI22_X1 U4193 ( .A1(n37809), .A2(n38788), .B1(n5474), .B2(n37181), .ZN(
        n6754) );
  OAI22_X1 U4194 ( .A1(n37809), .A2(n38795), .B1(n5474), .B2(n37182), .ZN(
        n6755) );
  OAI22_X1 U4195 ( .A1(n37809), .A2(n38802), .B1(n5474), .B2(n37183), .ZN(
        n6756) );
  OAI22_X1 U4196 ( .A1(n37809), .A2(n38809), .B1(n5474), .B2(n37184), .ZN(
        n6757) );
  OAI22_X1 U4197 ( .A1(n37809), .A2(n38816), .B1(n5474), .B2(n37185), .ZN(
        n6758) );
  OAI22_X1 U4198 ( .A1(n37810), .A2(n38823), .B1(n5474), .B2(n37186), .ZN(
        n6759) );
  OAI22_X1 U4199 ( .A1(n37810), .A2(n38830), .B1(n37805), .B2(n37187), .ZN(
        n6760) );
  OAI22_X1 U4200 ( .A1(n37810), .A2(n38837), .B1(n37805), .B2(n37188), .ZN(
        n6761) );
  OAI22_X1 U4201 ( .A1(n37810), .A2(n38844), .B1(n37805), .B2(n37189), .ZN(
        n6762) );
  OAI22_X1 U4202 ( .A1(n37851), .A2(n38683), .B1(n37850), .B2(n36782), .ZN(
        n6867) );
  OAI22_X1 U4203 ( .A1(n37851), .A2(n38690), .B1(n37850), .B2(n36783), .ZN(
        n6868) );
  OAI22_X1 U4204 ( .A1(n37851), .A2(n38697), .B1(n37850), .B2(n36784), .ZN(
        n6869) );
  OAI22_X1 U4205 ( .A1(n37851), .A2(n38704), .B1(n37850), .B2(n36785), .ZN(
        n6870) );
  OAI22_X1 U4206 ( .A1(n37851), .A2(n38711), .B1(n37850), .B2(n36786), .ZN(
        n6871) );
  OAI22_X1 U4207 ( .A1(n37852), .A2(n38718), .B1(n37850), .B2(n36787), .ZN(
        n6872) );
  OAI22_X1 U4208 ( .A1(n37852), .A2(n38725), .B1(n37850), .B2(n36788), .ZN(
        n6873) );
  OAI22_X1 U4209 ( .A1(n37852), .A2(n38732), .B1(n37850), .B2(n36789), .ZN(
        n6874) );
  OAI22_X1 U4210 ( .A1(n37852), .A2(n38739), .B1(n37850), .B2(n36790), .ZN(
        n6875) );
  OAI22_X1 U4211 ( .A1(n37852), .A2(n38746), .B1(n37850), .B2(n36791), .ZN(
        n6876) );
  OAI22_X1 U4212 ( .A1(n37853), .A2(n38753), .B1(n37850), .B2(n36792), .ZN(
        n6877) );
  OAI22_X1 U4213 ( .A1(n37853), .A2(n38760), .B1(n37850), .B2(n36793), .ZN(
        n6878) );
  OAI22_X1 U4214 ( .A1(n37853), .A2(n38767), .B1(n37850), .B2(n36794), .ZN(
        n6879) );
  OAI22_X1 U4215 ( .A1(n37853), .A2(n38774), .B1(n37850), .B2(n36795), .ZN(
        n6880) );
  OAI22_X1 U4216 ( .A1(n37853), .A2(n38781), .B1(n5334), .B2(n36796), .ZN(
        n6881) );
  OAI22_X1 U4217 ( .A1(n37854), .A2(n38788), .B1(n5334), .B2(n36797), .ZN(
        n6882) );
  OAI22_X1 U4218 ( .A1(n37854), .A2(n38795), .B1(n5334), .B2(n36798), .ZN(
        n6883) );
  OAI22_X1 U4219 ( .A1(n37854), .A2(n38802), .B1(n5334), .B2(n36799), .ZN(
        n6884) );
  OAI22_X1 U4220 ( .A1(n37854), .A2(n38809), .B1(n5334), .B2(n36800), .ZN(
        n6885) );
  OAI22_X1 U4221 ( .A1(n37854), .A2(n38816), .B1(n5334), .B2(n36801), .ZN(
        n6886) );
  OAI22_X1 U4222 ( .A1(n37855), .A2(n38823), .B1(n5334), .B2(n36802), .ZN(
        n6887) );
  OAI22_X1 U4223 ( .A1(n37855), .A2(n38830), .B1(n37850), .B2(n36803), .ZN(
        n6888) );
  OAI22_X1 U4224 ( .A1(n37855), .A2(n38837), .B1(n37850), .B2(n36804), .ZN(
        n6889) );
  OAI22_X1 U4225 ( .A1(n37855), .A2(n38844), .B1(n37850), .B2(n36805), .ZN(
        n6890) );
  OAI22_X1 U4226 ( .A1(n37860), .A2(n38683), .B1(n37859), .B2(n37190), .ZN(
        n6899) );
  OAI22_X1 U4227 ( .A1(n37860), .A2(n38690), .B1(n37859), .B2(n37191), .ZN(
        n6900) );
  OAI22_X1 U4228 ( .A1(n37860), .A2(n38697), .B1(n37859), .B2(n37192), .ZN(
        n6901) );
  OAI22_X1 U4229 ( .A1(n37860), .A2(n38704), .B1(n37859), .B2(n37193), .ZN(
        n6902) );
  OAI22_X1 U4230 ( .A1(n37860), .A2(n38711), .B1(n37859), .B2(n37194), .ZN(
        n6903) );
  OAI22_X1 U4231 ( .A1(n37861), .A2(n38718), .B1(n37859), .B2(n37195), .ZN(
        n6904) );
  OAI22_X1 U4232 ( .A1(n37861), .A2(n38725), .B1(n37859), .B2(n37196), .ZN(
        n6905) );
  OAI22_X1 U4233 ( .A1(n37861), .A2(n38732), .B1(n37859), .B2(n37197), .ZN(
        n6906) );
  OAI22_X1 U4234 ( .A1(n37861), .A2(n38739), .B1(n37859), .B2(n37198), .ZN(
        n6907) );
  OAI22_X1 U4235 ( .A1(n37861), .A2(n38746), .B1(n37859), .B2(n37199), .ZN(
        n6908) );
  OAI22_X1 U4236 ( .A1(n37862), .A2(n38753), .B1(n37859), .B2(n37200), .ZN(
        n6909) );
  OAI22_X1 U4237 ( .A1(n37862), .A2(n38760), .B1(n37859), .B2(n37201), .ZN(
        n6910) );
  OAI22_X1 U4238 ( .A1(n37862), .A2(n38767), .B1(n37859), .B2(n37202), .ZN(
        n6911) );
  OAI22_X1 U4239 ( .A1(n37862), .A2(n38774), .B1(n37859), .B2(n37203), .ZN(
        n6912) );
  OAI22_X1 U4240 ( .A1(n37862), .A2(n38781), .B1(n5299), .B2(n37204), .ZN(
        n6913) );
  OAI22_X1 U4241 ( .A1(n37863), .A2(n38788), .B1(n5299), .B2(n37205), .ZN(
        n6914) );
  OAI22_X1 U4242 ( .A1(n37863), .A2(n38795), .B1(n5299), .B2(n37206), .ZN(
        n6915) );
  OAI22_X1 U4243 ( .A1(n37863), .A2(n38802), .B1(n5299), .B2(n37207), .ZN(
        n6916) );
  OAI22_X1 U4244 ( .A1(n37863), .A2(n38809), .B1(n5299), .B2(n37208), .ZN(
        n6917) );
  OAI22_X1 U4245 ( .A1(n37863), .A2(n38816), .B1(n5299), .B2(n37209), .ZN(
        n6918) );
  OAI22_X1 U4246 ( .A1(n37864), .A2(n38823), .B1(n5299), .B2(n37210), .ZN(
        n6919) );
  OAI22_X1 U4247 ( .A1(n37864), .A2(n38830), .B1(n37859), .B2(n37211), .ZN(
        n6920) );
  OAI22_X1 U4248 ( .A1(n37864), .A2(n38837), .B1(n37859), .B2(n37212), .ZN(
        n6921) );
  OAI22_X1 U4249 ( .A1(n37864), .A2(n38844), .B1(n37859), .B2(n37213), .ZN(
        n6922) );
  OAI22_X1 U4250 ( .A1(n37905), .A2(n38683), .B1(n37904), .B2(n36806), .ZN(
        n7027) );
  OAI22_X1 U4251 ( .A1(n37905), .A2(n38690), .B1(n37904), .B2(n36807), .ZN(
        n7028) );
  OAI22_X1 U4252 ( .A1(n37905), .A2(n38697), .B1(n37904), .B2(n36808), .ZN(
        n7029) );
  OAI22_X1 U4253 ( .A1(n37905), .A2(n38704), .B1(n37904), .B2(n36809), .ZN(
        n7030) );
  OAI22_X1 U4254 ( .A1(n37905), .A2(n38711), .B1(n37904), .B2(n36810), .ZN(
        n7031) );
  OAI22_X1 U4255 ( .A1(n37906), .A2(n38718), .B1(n37904), .B2(n36811), .ZN(
        n7032) );
  OAI22_X1 U4256 ( .A1(n37906), .A2(n38725), .B1(n37904), .B2(n36812), .ZN(
        n7033) );
  OAI22_X1 U4257 ( .A1(n37906), .A2(n38732), .B1(n37904), .B2(n36813), .ZN(
        n7034) );
  OAI22_X1 U4258 ( .A1(n37906), .A2(n38739), .B1(n37904), .B2(n36814), .ZN(
        n7035) );
  OAI22_X1 U4259 ( .A1(n37906), .A2(n38746), .B1(n37904), .B2(n36815), .ZN(
        n7036) );
  OAI22_X1 U4260 ( .A1(n37907), .A2(n38753), .B1(n37904), .B2(n36816), .ZN(
        n7037) );
  OAI22_X1 U4261 ( .A1(n37907), .A2(n38760), .B1(n37904), .B2(n36817), .ZN(
        n7038) );
  OAI22_X1 U4262 ( .A1(n37907), .A2(n38767), .B1(n37904), .B2(n36818), .ZN(
        n7039) );
  OAI22_X1 U4263 ( .A1(n37907), .A2(n38774), .B1(n37904), .B2(n36819), .ZN(
        n7040) );
  OAI22_X1 U4264 ( .A1(n37907), .A2(n38781), .B1(n5159), .B2(n36820), .ZN(
        n7041) );
  OAI22_X1 U4265 ( .A1(n37908), .A2(n38788), .B1(n5159), .B2(n36821), .ZN(
        n7042) );
  OAI22_X1 U4266 ( .A1(n37908), .A2(n38795), .B1(n5159), .B2(n36822), .ZN(
        n7043) );
  OAI22_X1 U4267 ( .A1(n37908), .A2(n38802), .B1(n5159), .B2(n36823), .ZN(
        n7044) );
  OAI22_X1 U4268 ( .A1(n37908), .A2(n38809), .B1(n5159), .B2(n36824), .ZN(
        n7045) );
  OAI22_X1 U4269 ( .A1(n37908), .A2(n38816), .B1(n5159), .B2(n36825), .ZN(
        n7046) );
  OAI22_X1 U4270 ( .A1(n37909), .A2(n38823), .B1(n5159), .B2(n36826), .ZN(
        n7047) );
  OAI22_X1 U4271 ( .A1(n37909), .A2(n38830), .B1(n37904), .B2(n36827), .ZN(
        n7048) );
  OAI22_X1 U4272 ( .A1(n37909), .A2(n38837), .B1(n37904), .B2(n36828), .ZN(
        n7049) );
  OAI22_X1 U4273 ( .A1(n37909), .A2(n38844), .B1(n37904), .B2(n36829), .ZN(
        n7050) );
  OAI22_X1 U4274 ( .A1(n37914), .A2(n38683), .B1(n37913), .B2(n37214), .ZN(
        n7059) );
  OAI22_X1 U4275 ( .A1(n37914), .A2(n38690), .B1(n37913), .B2(n37215), .ZN(
        n7060) );
  OAI22_X1 U4276 ( .A1(n37914), .A2(n38697), .B1(n37913), .B2(n37216), .ZN(
        n7061) );
  OAI22_X1 U4277 ( .A1(n37914), .A2(n38704), .B1(n37913), .B2(n37217), .ZN(
        n7062) );
  OAI22_X1 U4278 ( .A1(n37914), .A2(n38711), .B1(n37913), .B2(n37218), .ZN(
        n7063) );
  OAI22_X1 U4279 ( .A1(n37915), .A2(n38718), .B1(n37913), .B2(n37219), .ZN(
        n7064) );
  OAI22_X1 U4280 ( .A1(n37915), .A2(n38725), .B1(n37913), .B2(n37220), .ZN(
        n7065) );
  OAI22_X1 U4281 ( .A1(n37915), .A2(n38732), .B1(n37913), .B2(n37221), .ZN(
        n7066) );
  OAI22_X1 U4282 ( .A1(n37915), .A2(n38739), .B1(n37913), .B2(n37222), .ZN(
        n7067) );
  OAI22_X1 U4283 ( .A1(n37915), .A2(n38746), .B1(n37913), .B2(n37223), .ZN(
        n7068) );
  OAI22_X1 U4284 ( .A1(n37916), .A2(n38753), .B1(n37913), .B2(n37224), .ZN(
        n7069) );
  OAI22_X1 U4285 ( .A1(n37916), .A2(n38760), .B1(n37913), .B2(n37225), .ZN(
        n7070) );
  OAI22_X1 U4286 ( .A1(n37916), .A2(n38767), .B1(n37913), .B2(n37226), .ZN(
        n7071) );
  OAI22_X1 U4287 ( .A1(n37916), .A2(n38774), .B1(n37913), .B2(n37227), .ZN(
        n7072) );
  OAI22_X1 U4288 ( .A1(n37916), .A2(n38781), .B1(n5124), .B2(n37228), .ZN(
        n7073) );
  OAI22_X1 U4289 ( .A1(n37917), .A2(n38788), .B1(n5124), .B2(n37229), .ZN(
        n7074) );
  OAI22_X1 U4290 ( .A1(n37917), .A2(n38795), .B1(n5124), .B2(n37230), .ZN(
        n7075) );
  OAI22_X1 U4291 ( .A1(n37917), .A2(n38802), .B1(n5124), .B2(n37231), .ZN(
        n7076) );
  OAI22_X1 U4292 ( .A1(n37917), .A2(n38809), .B1(n5124), .B2(n37232), .ZN(
        n7077) );
  OAI22_X1 U4293 ( .A1(n37917), .A2(n38816), .B1(n5124), .B2(n37233), .ZN(
        n7078) );
  OAI22_X1 U4294 ( .A1(n37918), .A2(n38823), .B1(n5124), .B2(n37234), .ZN(
        n7079) );
  OAI22_X1 U4295 ( .A1(n37918), .A2(n38830), .B1(n37913), .B2(n37235), .ZN(
        n7080) );
  OAI22_X1 U4296 ( .A1(n37918), .A2(n38837), .B1(n37913), .B2(n37236), .ZN(
        n7081) );
  OAI22_X1 U4297 ( .A1(n37918), .A2(n38844), .B1(n37913), .B2(n37237), .ZN(
        n7082) );
  OAI22_X1 U4298 ( .A1(n37959), .A2(n38682), .B1(n37958), .B2(n36830), .ZN(
        n7187) );
  OAI22_X1 U4299 ( .A1(n37959), .A2(n38689), .B1(n37958), .B2(n36831), .ZN(
        n7188) );
  OAI22_X1 U4300 ( .A1(n37959), .A2(n38696), .B1(n37958), .B2(n36832), .ZN(
        n7189) );
  OAI22_X1 U4301 ( .A1(n37959), .A2(n38703), .B1(n37958), .B2(n36833), .ZN(
        n7190) );
  OAI22_X1 U4302 ( .A1(n37959), .A2(n38710), .B1(n37958), .B2(n36834), .ZN(
        n7191) );
  OAI22_X1 U4303 ( .A1(n37960), .A2(n38717), .B1(n37958), .B2(n36835), .ZN(
        n7192) );
  OAI22_X1 U4304 ( .A1(n37960), .A2(n38724), .B1(n37958), .B2(n36836), .ZN(
        n7193) );
  OAI22_X1 U4305 ( .A1(n37960), .A2(n38731), .B1(n37958), .B2(n36837), .ZN(
        n7194) );
  OAI22_X1 U4306 ( .A1(n37960), .A2(n38738), .B1(n37958), .B2(n36838), .ZN(
        n7195) );
  OAI22_X1 U4307 ( .A1(n37960), .A2(n38745), .B1(n37958), .B2(n36839), .ZN(
        n7196) );
  OAI22_X1 U4308 ( .A1(n37961), .A2(n38752), .B1(n37958), .B2(n36840), .ZN(
        n7197) );
  OAI22_X1 U4309 ( .A1(n37961), .A2(n38759), .B1(n37958), .B2(n36841), .ZN(
        n7198) );
  OAI22_X1 U4310 ( .A1(n37961), .A2(n38766), .B1(n37958), .B2(n36842), .ZN(
        n7199) );
  OAI22_X1 U4311 ( .A1(n37961), .A2(n38773), .B1(n37958), .B2(n36843), .ZN(
        n7200) );
  OAI22_X1 U4312 ( .A1(n37961), .A2(n38780), .B1(n4983), .B2(n36844), .ZN(
        n7201) );
  OAI22_X1 U4313 ( .A1(n37962), .A2(n38787), .B1(n4983), .B2(n36845), .ZN(
        n7202) );
  OAI22_X1 U4314 ( .A1(n37962), .A2(n38794), .B1(n4983), .B2(n36846), .ZN(
        n7203) );
  OAI22_X1 U4315 ( .A1(n37962), .A2(n38801), .B1(n4983), .B2(n36847), .ZN(
        n7204) );
  OAI22_X1 U4316 ( .A1(n37962), .A2(n38808), .B1(n4983), .B2(n36848), .ZN(
        n7205) );
  OAI22_X1 U4317 ( .A1(n37962), .A2(n38815), .B1(n4983), .B2(n36849), .ZN(
        n7206) );
  OAI22_X1 U4318 ( .A1(n37963), .A2(n38822), .B1(n4983), .B2(n36850), .ZN(
        n7207) );
  OAI22_X1 U4319 ( .A1(n37963), .A2(n38829), .B1(n37958), .B2(n36851), .ZN(
        n7208) );
  OAI22_X1 U4320 ( .A1(n37963), .A2(n38836), .B1(n37958), .B2(n36852), .ZN(
        n7209) );
  OAI22_X1 U4321 ( .A1(n37963), .A2(n38843), .B1(n37958), .B2(n36853), .ZN(
        n7210) );
  OAI22_X1 U4322 ( .A1(n37992), .A2(n38682), .B1(n37991), .B2(n36854), .ZN(
        n7283) );
  OAI22_X1 U4323 ( .A1(n37992), .A2(n38689), .B1(n37991), .B2(n36855), .ZN(
        n7284) );
  OAI22_X1 U4324 ( .A1(n37992), .A2(n38696), .B1(n37991), .B2(n36856), .ZN(
        n7285) );
  OAI22_X1 U4325 ( .A1(n37992), .A2(n38703), .B1(n37991), .B2(n36857), .ZN(
        n7286) );
  OAI22_X1 U4326 ( .A1(n37992), .A2(n38710), .B1(n37991), .B2(n36858), .ZN(
        n7287) );
  OAI22_X1 U4327 ( .A1(n37993), .A2(n38717), .B1(n37991), .B2(n36859), .ZN(
        n7288) );
  OAI22_X1 U4328 ( .A1(n37993), .A2(n38724), .B1(n37991), .B2(n36860), .ZN(
        n7289) );
  OAI22_X1 U4329 ( .A1(n37993), .A2(n38731), .B1(n37991), .B2(n36861), .ZN(
        n7290) );
  OAI22_X1 U4330 ( .A1(n37993), .A2(n38738), .B1(n37991), .B2(n36862), .ZN(
        n7291) );
  OAI22_X1 U4331 ( .A1(n37993), .A2(n38745), .B1(n37991), .B2(n36863), .ZN(
        n7292) );
  OAI22_X1 U4332 ( .A1(n37994), .A2(n38752), .B1(n37991), .B2(n36864), .ZN(
        n7293) );
  OAI22_X1 U4333 ( .A1(n37994), .A2(n38759), .B1(n37991), .B2(n36865), .ZN(
        n7294) );
  OAI22_X1 U4334 ( .A1(n37994), .A2(n38766), .B1(n37991), .B2(n36866), .ZN(
        n7295) );
  OAI22_X1 U4335 ( .A1(n37994), .A2(n38773), .B1(n37991), .B2(n36867), .ZN(
        n7296) );
  OAI22_X1 U4336 ( .A1(n37994), .A2(n38780), .B1(n4878), .B2(n36868), .ZN(
        n7297) );
  OAI22_X1 U4337 ( .A1(n37995), .A2(n38787), .B1(n4878), .B2(n36869), .ZN(
        n7298) );
  OAI22_X1 U4338 ( .A1(n37995), .A2(n38794), .B1(n4878), .B2(n36870), .ZN(
        n7299) );
  OAI22_X1 U4339 ( .A1(n37995), .A2(n38801), .B1(n4878), .B2(n36871), .ZN(
        n7300) );
  OAI22_X1 U4340 ( .A1(n37995), .A2(n38808), .B1(n4878), .B2(n36872), .ZN(
        n7301) );
  OAI22_X1 U4341 ( .A1(n37995), .A2(n38815), .B1(n4878), .B2(n36873), .ZN(
        n7302) );
  OAI22_X1 U4342 ( .A1(n37996), .A2(n38822), .B1(n4878), .B2(n36874), .ZN(
        n7303) );
  OAI22_X1 U4343 ( .A1(n37996), .A2(n38829), .B1(n37991), .B2(n36875), .ZN(
        n7304) );
  OAI22_X1 U4344 ( .A1(n37996), .A2(n38836), .B1(n37991), .B2(n36876), .ZN(
        n7305) );
  OAI22_X1 U4345 ( .A1(n37996), .A2(n38843), .B1(n37991), .B2(n36877), .ZN(
        n7306) );
  OAI22_X1 U4346 ( .A1(n38013), .A2(n38681), .B1(n38012), .B2(n37238), .ZN(
        n7347) );
  OAI22_X1 U4347 ( .A1(n38013), .A2(n38688), .B1(n38012), .B2(n37239), .ZN(
        n7348) );
  OAI22_X1 U4348 ( .A1(n38013), .A2(n38695), .B1(n38012), .B2(n37240), .ZN(
        n7349) );
  OAI22_X1 U4349 ( .A1(n38013), .A2(n38702), .B1(n38012), .B2(n37241), .ZN(
        n7350) );
  OAI22_X1 U4350 ( .A1(n38013), .A2(n38709), .B1(n38012), .B2(n37242), .ZN(
        n7351) );
  OAI22_X1 U4351 ( .A1(n38014), .A2(n38716), .B1(n38012), .B2(n37243), .ZN(
        n7352) );
  OAI22_X1 U4352 ( .A1(n38014), .A2(n38723), .B1(n38012), .B2(n37244), .ZN(
        n7353) );
  OAI22_X1 U4353 ( .A1(n38014), .A2(n38730), .B1(n38012), .B2(n37245), .ZN(
        n7354) );
  OAI22_X1 U4354 ( .A1(n38014), .A2(n38737), .B1(n38012), .B2(n37246), .ZN(
        n7355) );
  OAI22_X1 U4355 ( .A1(n38014), .A2(n38744), .B1(n38012), .B2(n37247), .ZN(
        n7356) );
  OAI22_X1 U4356 ( .A1(n38015), .A2(n38751), .B1(n38012), .B2(n37248), .ZN(
        n7357) );
  OAI22_X1 U4357 ( .A1(n38015), .A2(n38758), .B1(n38012), .B2(n37249), .ZN(
        n7358) );
  OAI22_X1 U4358 ( .A1(n38015), .A2(n38765), .B1(n38012), .B2(n37250), .ZN(
        n7359) );
  OAI22_X1 U4359 ( .A1(n38015), .A2(n38772), .B1(n38012), .B2(n37251), .ZN(
        n7360) );
  OAI22_X1 U4360 ( .A1(n38015), .A2(n38779), .B1(n4808), .B2(n37252), .ZN(
        n7361) );
  OAI22_X1 U4361 ( .A1(n38016), .A2(n38786), .B1(n4808), .B2(n37253), .ZN(
        n7362) );
  OAI22_X1 U4362 ( .A1(n38016), .A2(n38793), .B1(n4808), .B2(n37254), .ZN(
        n7363) );
  OAI22_X1 U4363 ( .A1(n38016), .A2(n38800), .B1(n4808), .B2(n37255), .ZN(
        n7364) );
  OAI22_X1 U4364 ( .A1(n38016), .A2(n38807), .B1(n4808), .B2(n37256), .ZN(
        n7365) );
  OAI22_X1 U4365 ( .A1(n38016), .A2(n38814), .B1(n4808), .B2(n37257), .ZN(
        n7366) );
  OAI22_X1 U4366 ( .A1(n38017), .A2(n38821), .B1(n4808), .B2(n37258), .ZN(
        n7367) );
  OAI22_X1 U4367 ( .A1(n38017), .A2(n38828), .B1(n38012), .B2(n37259), .ZN(
        n7368) );
  OAI22_X1 U4368 ( .A1(n38017), .A2(n38835), .B1(n38012), .B2(n37260), .ZN(
        n7369) );
  OAI22_X1 U4369 ( .A1(n38017), .A2(n38842), .B1(n38012), .B2(n37261), .ZN(
        n7370) );
  OAI22_X1 U4370 ( .A1(n38046), .A2(n38682), .B1(n38045), .B2(n36878), .ZN(
        n7443) );
  OAI22_X1 U4371 ( .A1(n38046), .A2(n38689), .B1(n38045), .B2(n36879), .ZN(
        n7444) );
  OAI22_X1 U4372 ( .A1(n38046), .A2(n38696), .B1(n38045), .B2(n36880), .ZN(
        n7445) );
  OAI22_X1 U4373 ( .A1(n38046), .A2(n38703), .B1(n38045), .B2(n36881), .ZN(
        n7446) );
  OAI22_X1 U4374 ( .A1(n38046), .A2(n38710), .B1(n38045), .B2(n36882), .ZN(
        n7447) );
  OAI22_X1 U4375 ( .A1(n38047), .A2(n38717), .B1(n38045), .B2(n36883), .ZN(
        n7448) );
  OAI22_X1 U4376 ( .A1(n38047), .A2(n38724), .B1(n38045), .B2(n36884), .ZN(
        n7449) );
  OAI22_X1 U4377 ( .A1(n38047), .A2(n38731), .B1(n38045), .B2(n36885), .ZN(
        n7450) );
  OAI22_X1 U4378 ( .A1(n38047), .A2(n38738), .B1(n38045), .B2(n36886), .ZN(
        n7451) );
  OAI22_X1 U4379 ( .A1(n38047), .A2(n38745), .B1(n38045), .B2(n36887), .ZN(
        n7452) );
  OAI22_X1 U4380 ( .A1(n38048), .A2(n38752), .B1(n38045), .B2(n36888), .ZN(
        n7453) );
  OAI22_X1 U4381 ( .A1(n38048), .A2(n38759), .B1(n38045), .B2(n36889), .ZN(
        n7454) );
  OAI22_X1 U4382 ( .A1(n38048), .A2(n38766), .B1(n38045), .B2(n36890), .ZN(
        n7455) );
  OAI22_X1 U4383 ( .A1(n38048), .A2(n38773), .B1(n38045), .B2(n36891), .ZN(
        n7456) );
  OAI22_X1 U4384 ( .A1(n38048), .A2(n38780), .B1(n4703), .B2(n36892), .ZN(
        n7457) );
  OAI22_X1 U4385 ( .A1(n38049), .A2(n38787), .B1(n4703), .B2(n36893), .ZN(
        n7458) );
  OAI22_X1 U4386 ( .A1(n38049), .A2(n38794), .B1(n4703), .B2(n36894), .ZN(
        n7459) );
  OAI22_X1 U4387 ( .A1(n38049), .A2(n38801), .B1(n4703), .B2(n36895), .ZN(
        n7460) );
  OAI22_X1 U4388 ( .A1(n38049), .A2(n38808), .B1(n4703), .B2(n36896), .ZN(
        n7461) );
  OAI22_X1 U4389 ( .A1(n38049), .A2(n38815), .B1(n4703), .B2(n36897), .ZN(
        n7462) );
  OAI22_X1 U4390 ( .A1(n38050), .A2(n38822), .B1(n4703), .B2(n36898), .ZN(
        n7463) );
  OAI22_X1 U4391 ( .A1(n38050), .A2(n38829), .B1(n38045), .B2(n36899), .ZN(
        n7464) );
  OAI22_X1 U4392 ( .A1(n38050), .A2(n38836), .B1(n38045), .B2(n36900), .ZN(
        n7465) );
  OAI22_X1 U4393 ( .A1(n38050), .A2(n38843), .B1(n38045), .B2(n36901), .ZN(
        n7466) );
  OAI22_X1 U4394 ( .A1(n38067), .A2(n38682), .B1(n38066), .B2(n37262), .ZN(
        n7507) );
  OAI22_X1 U4395 ( .A1(n38067), .A2(n38689), .B1(n38066), .B2(n37263), .ZN(
        n7508) );
  OAI22_X1 U4396 ( .A1(n38067), .A2(n38696), .B1(n38066), .B2(n37264), .ZN(
        n7509) );
  OAI22_X1 U4397 ( .A1(n38067), .A2(n38703), .B1(n38066), .B2(n37265), .ZN(
        n7510) );
  OAI22_X1 U4398 ( .A1(n38067), .A2(n38710), .B1(n38066), .B2(n37266), .ZN(
        n7511) );
  OAI22_X1 U4399 ( .A1(n38068), .A2(n38717), .B1(n38066), .B2(n37267), .ZN(
        n7512) );
  OAI22_X1 U4400 ( .A1(n38068), .A2(n38724), .B1(n38066), .B2(n37268), .ZN(
        n7513) );
  OAI22_X1 U4401 ( .A1(n38068), .A2(n38731), .B1(n38066), .B2(n37269), .ZN(
        n7514) );
  OAI22_X1 U4402 ( .A1(n38068), .A2(n38738), .B1(n38066), .B2(n37270), .ZN(
        n7515) );
  OAI22_X1 U4403 ( .A1(n38068), .A2(n38745), .B1(n38066), .B2(n37271), .ZN(
        n7516) );
  OAI22_X1 U4404 ( .A1(n38069), .A2(n38752), .B1(n38066), .B2(n37272), .ZN(
        n7517) );
  OAI22_X1 U4405 ( .A1(n38069), .A2(n38759), .B1(n38066), .B2(n37273), .ZN(
        n7518) );
  OAI22_X1 U4406 ( .A1(n38069), .A2(n38766), .B1(n38066), .B2(n37274), .ZN(
        n7519) );
  OAI22_X1 U4407 ( .A1(n38069), .A2(n38773), .B1(n38066), .B2(n37275), .ZN(
        n7520) );
  OAI22_X1 U4408 ( .A1(n38069), .A2(n38780), .B1(n4633), .B2(n37276), .ZN(
        n7521) );
  OAI22_X1 U4409 ( .A1(n38070), .A2(n38787), .B1(n4633), .B2(n37277), .ZN(
        n7522) );
  OAI22_X1 U4410 ( .A1(n38070), .A2(n38794), .B1(n4633), .B2(n37278), .ZN(
        n7523) );
  OAI22_X1 U4411 ( .A1(n38070), .A2(n38801), .B1(n4633), .B2(n37279), .ZN(
        n7524) );
  OAI22_X1 U4412 ( .A1(n38070), .A2(n38808), .B1(n4633), .B2(n37280), .ZN(
        n7525) );
  OAI22_X1 U4413 ( .A1(n38070), .A2(n38815), .B1(n4633), .B2(n37281), .ZN(
        n7526) );
  OAI22_X1 U4414 ( .A1(n38071), .A2(n38822), .B1(n4633), .B2(n37282), .ZN(
        n7527) );
  OAI22_X1 U4415 ( .A1(n38071), .A2(n38829), .B1(n38066), .B2(n37283), .ZN(
        n7528) );
  OAI22_X1 U4416 ( .A1(n38071), .A2(n38836), .B1(n38066), .B2(n37284), .ZN(
        n7529) );
  OAI22_X1 U4417 ( .A1(n38071), .A2(n38843), .B1(n38066), .B2(n37285), .ZN(
        n7530) );
  OAI22_X1 U4418 ( .A1(n38100), .A2(n38681), .B1(n38099), .B2(n36902), .ZN(
        n7603) );
  OAI22_X1 U4419 ( .A1(n38100), .A2(n38688), .B1(n38099), .B2(n36903), .ZN(
        n7604) );
  OAI22_X1 U4420 ( .A1(n38100), .A2(n38695), .B1(n38099), .B2(n36904), .ZN(
        n7605) );
  OAI22_X1 U4421 ( .A1(n38100), .A2(n38702), .B1(n38099), .B2(n36905), .ZN(
        n7606) );
  OAI22_X1 U4422 ( .A1(n38100), .A2(n38709), .B1(n38099), .B2(n36906), .ZN(
        n7607) );
  OAI22_X1 U4423 ( .A1(n38101), .A2(n38716), .B1(n38099), .B2(n36907), .ZN(
        n7608) );
  OAI22_X1 U4424 ( .A1(n38101), .A2(n38723), .B1(n38099), .B2(n36908), .ZN(
        n7609) );
  OAI22_X1 U4425 ( .A1(n38101), .A2(n38730), .B1(n38099), .B2(n36909), .ZN(
        n7610) );
  OAI22_X1 U4426 ( .A1(n38101), .A2(n38737), .B1(n38099), .B2(n36910), .ZN(
        n7611) );
  OAI22_X1 U4427 ( .A1(n38101), .A2(n38744), .B1(n38099), .B2(n36911), .ZN(
        n7612) );
  OAI22_X1 U4428 ( .A1(n38102), .A2(n38751), .B1(n38099), .B2(n36912), .ZN(
        n7613) );
  OAI22_X1 U4429 ( .A1(n38102), .A2(n38758), .B1(n38099), .B2(n36913), .ZN(
        n7614) );
  OAI22_X1 U4430 ( .A1(n38102), .A2(n38765), .B1(n38099), .B2(n36914), .ZN(
        n7615) );
  OAI22_X1 U4431 ( .A1(n38102), .A2(n38772), .B1(n38099), .B2(n36915), .ZN(
        n7616) );
  OAI22_X1 U4432 ( .A1(n38102), .A2(n38779), .B1(n4528), .B2(n36916), .ZN(
        n7617) );
  OAI22_X1 U4433 ( .A1(n38103), .A2(n38786), .B1(n4528), .B2(n36917), .ZN(
        n7618) );
  OAI22_X1 U4434 ( .A1(n38103), .A2(n38793), .B1(n4528), .B2(n36918), .ZN(
        n7619) );
  OAI22_X1 U4435 ( .A1(n38103), .A2(n38800), .B1(n4528), .B2(n36919), .ZN(
        n7620) );
  OAI22_X1 U4436 ( .A1(n38103), .A2(n38807), .B1(n4528), .B2(n36920), .ZN(
        n7621) );
  OAI22_X1 U4437 ( .A1(n38103), .A2(n38814), .B1(n4528), .B2(n36921), .ZN(
        n7622) );
  OAI22_X1 U4438 ( .A1(n38104), .A2(n38821), .B1(n4528), .B2(n36922), .ZN(
        n7623) );
  OAI22_X1 U4439 ( .A1(n38104), .A2(n38828), .B1(n38099), .B2(n36923), .ZN(
        n7624) );
  OAI22_X1 U4440 ( .A1(n38104), .A2(n38835), .B1(n38099), .B2(n36924), .ZN(
        n7625) );
  OAI22_X1 U4441 ( .A1(n38104), .A2(n38842), .B1(n38099), .B2(n36925), .ZN(
        n7626) );
  OAI22_X1 U4442 ( .A1(n38121), .A2(n38681), .B1(n38120), .B2(n37286), .ZN(
        n7667) );
  OAI22_X1 U4443 ( .A1(n38121), .A2(n38688), .B1(n38120), .B2(n37287), .ZN(
        n7668) );
  OAI22_X1 U4444 ( .A1(n38121), .A2(n38695), .B1(n38120), .B2(n37288), .ZN(
        n7669) );
  OAI22_X1 U4445 ( .A1(n38121), .A2(n38702), .B1(n38120), .B2(n37289), .ZN(
        n7670) );
  OAI22_X1 U4446 ( .A1(n38121), .A2(n38709), .B1(n38120), .B2(n37290), .ZN(
        n7671) );
  OAI22_X1 U4447 ( .A1(n38122), .A2(n38716), .B1(n38120), .B2(n37291), .ZN(
        n7672) );
  OAI22_X1 U4448 ( .A1(n38122), .A2(n38723), .B1(n38120), .B2(n37292), .ZN(
        n7673) );
  OAI22_X1 U4449 ( .A1(n38122), .A2(n38730), .B1(n38120), .B2(n37293), .ZN(
        n7674) );
  OAI22_X1 U4450 ( .A1(n38122), .A2(n38737), .B1(n38120), .B2(n37294), .ZN(
        n7675) );
  OAI22_X1 U4451 ( .A1(n38122), .A2(n38744), .B1(n38120), .B2(n37295), .ZN(
        n7676) );
  OAI22_X1 U4452 ( .A1(n38123), .A2(n38751), .B1(n38120), .B2(n37296), .ZN(
        n7677) );
  OAI22_X1 U4453 ( .A1(n38123), .A2(n38758), .B1(n38120), .B2(n37297), .ZN(
        n7678) );
  OAI22_X1 U4454 ( .A1(n38123), .A2(n38765), .B1(n38120), .B2(n37298), .ZN(
        n7679) );
  OAI22_X1 U4455 ( .A1(n38123), .A2(n38772), .B1(n38120), .B2(n37299), .ZN(
        n7680) );
  OAI22_X1 U4456 ( .A1(n38123), .A2(n38779), .B1(n4458), .B2(n37300), .ZN(
        n7681) );
  OAI22_X1 U4457 ( .A1(n38124), .A2(n38786), .B1(n4458), .B2(n37301), .ZN(
        n7682) );
  OAI22_X1 U4458 ( .A1(n38124), .A2(n38793), .B1(n4458), .B2(n37302), .ZN(
        n7683) );
  OAI22_X1 U4459 ( .A1(n38124), .A2(n38800), .B1(n4458), .B2(n37303), .ZN(
        n7684) );
  OAI22_X1 U4460 ( .A1(n38124), .A2(n38807), .B1(n4458), .B2(n37304), .ZN(
        n7685) );
  OAI22_X1 U4461 ( .A1(n38124), .A2(n38814), .B1(n4458), .B2(n37305), .ZN(
        n7686) );
  OAI22_X1 U4462 ( .A1(n38125), .A2(n38821), .B1(n4458), .B2(n37306), .ZN(
        n7687) );
  OAI22_X1 U4463 ( .A1(n38125), .A2(n38828), .B1(n38120), .B2(n37307), .ZN(
        n7688) );
  OAI22_X1 U4464 ( .A1(n38125), .A2(n38835), .B1(n38120), .B2(n37308), .ZN(
        n7689) );
  OAI22_X1 U4465 ( .A1(n38125), .A2(n38842), .B1(n38120), .B2(n37309), .ZN(
        n7690) );
  OAI22_X1 U4466 ( .A1(n38154), .A2(n38681), .B1(n38153), .B2(n37310), .ZN(
        n7763) );
  OAI22_X1 U4467 ( .A1(n38154), .A2(n38688), .B1(n38153), .B2(n37311), .ZN(
        n7764) );
  OAI22_X1 U4468 ( .A1(n38154), .A2(n38695), .B1(n38153), .B2(n37312), .ZN(
        n7765) );
  OAI22_X1 U4469 ( .A1(n38154), .A2(n38702), .B1(n38153), .B2(n37313), .ZN(
        n7766) );
  OAI22_X1 U4470 ( .A1(n38154), .A2(n38709), .B1(n38153), .B2(n37314), .ZN(
        n7767) );
  OAI22_X1 U4471 ( .A1(n38155), .A2(n38716), .B1(n38153), .B2(n37315), .ZN(
        n7768) );
  OAI22_X1 U4472 ( .A1(n38155), .A2(n38723), .B1(n38153), .B2(n37316), .ZN(
        n7769) );
  OAI22_X1 U4473 ( .A1(n38155), .A2(n38730), .B1(n38153), .B2(n37317), .ZN(
        n7770) );
  OAI22_X1 U4474 ( .A1(n38155), .A2(n38737), .B1(n38153), .B2(n37318), .ZN(
        n7771) );
  OAI22_X1 U4475 ( .A1(n38155), .A2(n38744), .B1(n38153), .B2(n37319), .ZN(
        n7772) );
  OAI22_X1 U4476 ( .A1(n38156), .A2(n38751), .B1(n38153), .B2(n37320), .ZN(
        n7773) );
  OAI22_X1 U4477 ( .A1(n38156), .A2(n38758), .B1(n38153), .B2(n37321), .ZN(
        n7774) );
  OAI22_X1 U4478 ( .A1(n38156), .A2(n38765), .B1(n38153), .B2(n37322), .ZN(
        n7775) );
  OAI22_X1 U4479 ( .A1(n38156), .A2(n38772), .B1(n38153), .B2(n37323), .ZN(
        n7776) );
  OAI22_X1 U4480 ( .A1(n38156), .A2(n38779), .B1(n4353), .B2(n37324), .ZN(
        n7777) );
  OAI22_X1 U4481 ( .A1(n38157), .A2(n38786), .B1(n4353), .B2(n37325), .ZN(
        n7778) );
  OAI22_X1 U4482 ( .A1(n38157), .A2(n38793), .B1(n4353), .B2(n37326), .ZN(
        n7779) );
  OAI22_X1 U4483 ( .A1(n38157), .A2(n38800), .B1(n4353), .B2(n37327), .ZN(
        n7780) );
  OAI22_X1 U4484 ( .A1(n38157), .A2(n38807), .B1(n4353), .B2(n37328), .ZN(
        n7781) );
  OAI22_X1 U4485 ( .A1(n38157), .A2(n38814), .B1(n4353), .B2(n37329), .ZN(
        n7782) );
  OAI22_X1 U4486 ( .A1(n38158), .A2(n38821), .B1(n4353), .B2(n37330), .ZN(
        n7783) );
  OAI22_X1 U4487 ( .A1(n38158), .A2(n38828), .B1(n38153), .B2(n37331), .ZN(
        n7784) );
  OAI22_X1 U4488 ( .A1(n38158), .A2(n38835), .B1(n38153), .B2(n37332), .ZN(
        n7785) );
  OAI22_X1 U4489 ( .A1(n38158), .A2(n38842), .B1(n38153), .B2(n37333), .ZN(
        n7786) );
  OAI22_X1 U4490 ( .A1(n38187), .A2(n38681), .B1(n38186), .B2(n36926), .ZN(
        n7859) );
  OAI22_X1 U4491 ( .A1(n38187), .A2(n38688), .B1(n38186), .B2(n36927), .ZN(
        n7860) );
  OAI22_X1 U4492 ( .A1(n38187), .A2(n38695), .B1(n38186), .B2(n36928), .ZN(
        n7861) );
  OAI22_X1 U4493 ( .A1(n38187), .A2(n38702), .B1(n38186), .B2(n36929), .ZN(
        n7862) );
  OAI22_X1 U4494 ( .A1(n38187), .A2(n38709), .B1(n38186), .B2(n36930), .ZN(
        n7863) );
  OAI22_X1 U4495 ( .A1(n38188), .A2(n38716), .B1(n38186), .B2(n36931), .ZN(
        n7864) );
  OAI22_X1 U4496 ( .A1(n38188), .A2(n38723), .B1(n38186), .B2(n36932), .ZN(
        n7865) );
  OAI22_X1 U4497 ( .A1(n38188), .A2(n38730), .B1(n38186), .B2(n36933), .ZN(
        n7866) );
  OAI22_X1 U4498 ( .A1(n38188), .A2(n38737), .B1(n38186), .B2(n36934), .ZN(
        n7867) );
  OAI22_X1 U4499 ( .A1(n38188), .A2(n38744), .B1(n38186), .B2(n36935), .ZN(
        n7868) );
  OAI22_X1 U4500 ( .A1(n38189), .A2(n38751), .B1(n38186), .B2(n36936), .ZN(
        n7869) );
  OAI22_X1 U4501 ( .A1(n38189), .A2(n38758), .B1(n38186), .B2(n36937), .ZN(
        n7870) );
  OAI22_X1 U4502 ( .A1(n38189), .A2(n38765), .B1(n38186), .B2(n36938), .ZN(
        n7871) );
  OAI22_X1 U4503 ( .A1(n38189), .A2(n38772), .B1(n38186), .B2(n36939), .ZN(
        n7872) );
  OAI22_X1 U4504 ( .A1(n38189), .A2(n38779), .B1(n4248), .B2(n36940), .ZN(
        n7873) );
  OAI22_X1 U4505 ( .A1(n38190), .A2(n38786), .B1(n4248), .B2(n36941), .ZN(
        n7874) );
  OAI22_X1 U4506 ( .A1(n38190), .A2(n38793), .B1(n4248), .B2(n36942), .ZN(
        n7875) );
  OAI22_X1 U4507 ( .A1(n38190), .A2(n38800), .B1(n4248), .B2(n36943), .ZN(
        n7876) );
  OAI22_X1 U4508 ( .A1(n38190), .A2(n38807), .B1(n4248), .B2(n36944), .ZN(
        n7877) );
  OAI22_X1 U4509 ( .A1(n38190), .A2(n38814), .B1(n4248), .B2(n36945), .ZN(
        n7878) );
  OAI22_X1 U4510 ( .A1(n38191), .A2(n38821), .B1(n4248), .B2(n36946), .ZN(
        n7879) );
  OAI22_X1 U4511 ( .A1(n38191), .A2(n38828), .B1(n38186), .B2(n36947), .ZN(
        n7880) );
  OAI22_X1 U4512 ( .A1(n38191), .A2(n38835), .B1(n38186), .B2(n36948), .ZN(
        n7881) );
  OAI22_X1 U4513 ( .A1(n38191), .A2(n38842), .B1(n38186), .B2(n36949), .ZN(
        n7882) );
  OAI22_X1 U4514 ( .A1(n38208), .A2(n38680), .B1(n38207), .B2(n37334), .ZN(
        n7923) );
  OAI22_X1 U4515 ( .A1(n38208), .A2(n38687), .B1(n38207), .B2(n37335), .ZN(
        n7924) );
  OAI22_X1 U4516 ( .A1(n38208), .A2(n38694), .B1(n38207), .B2(n37336), .ZN(
        n7925) );
  OAI22_X1 U4517 ( .A1(n38208), .A2(n38701), .B1(n38207), .B2(n37337), .ZN(
        n7926) );
  OAI22_X1 U4518 ( .A1(n38208), .A2(n38708), .B1(n38207), .B2(n37338), .ZN(
        n7927) );
  OAI22_X1 U4519 ( .A1(n38209), .A2(n38715), .B1(n38207), .B2(n37339), .ZN(
        n7928) );
  OAI22_X1 U4520 ( .A1(n38209), .A2(n38722), .B1(n38207), .B2(n37340), .ZN(
        n7929) );
  OAI22_X1 U4521 ( .A1(n38209), .A2(n38729), .B1(n38207), .B2(n37341), .ZN(
        n7930) );
  OAI22_X1 U4522 ( .A1(n38209), .A2(n38736), .B1(n38207), .B2(n37342), .ZN(
        n7931) );
  OAI22_X1 U4523 ( .A1(n38209), .A2(n38743), .B1(n38207), .B2(n37343), .ZN(
        n7932) );
  OAI22_X1 U4524 ( .A1(n38210), .A2(n38750), .B1(n38207), .B2(n37344), .ZN(
        n7933) );
  OAI22_X1 U4525 ( .A1(n38210), .A2(n38757), .B1(n38207), .B2(n37345), .ZN(
        n7934) );
  OAI22_X1 U4526 ( .A1(n38210), .A2(n38764), .B1(n38207), .B2(n37346), .ZN(
        n7935) );
  OAI22_X1 U4527 ( .A1(n38210), .A2(n38771), .B1(n38207), .B2(n37347), .ZN(
        n7936) );
  OAI22_X1 U4528 ( .A1(n38210), .A2(n38778), .B1(n4178), .B2(n37348), .ZN(
        n7937) );
  OAI22_X1 U4529 ( .A1(n38211), .A2(n38785), .B1(n4178), .B2(n37349), .ZN(
        n7938) );
  OAI22_X1 U4530 ( .A1(n38211), .A2(n38792), .B1(n4178), .B2(n37350), .ZN(
        n7939) );
  OAI22_X1 U4531 ( .A1(n38211), .A2(n38799), .B1(n4178), .B2(n37351), .ZN(
        n7940) );
  OAI22_X1 U4532 ( .A1(n38211), .A2(n38806), .B1(n4178), .B2(n37352), .ZN(
        n7941) );
  OAI22_X1 U4533 ( .A1(n38211), .A2(n38813), .B1(n4178), .B2(n37353), .ZN(
        n7942) );
  OAI22_X1 U4534 ( .A1(n38212), .A2(n38820), .B1(n4178), .B2(n37354), .ZN(
        n7943) );
  OAI22_X1 U4535 ( .A1(n38212), .A2(n38827), .B1(n38207), .B2(n37355), .ZN(
        n7944) );
  OAI22_X1 U4536 ( .A1(n38212), .A2(n38834), .B1(n38207), .B2(n37356), .ZN(
        n7945) );
  OAI22_X1 U4537 ( .A1(n38212), .A2(n38841), .B1(n38207), .B2(n37357), .ZN(
        n7946) );
  OAI22_X1 U4538 ( .A1(n38241), .A2(n38680), .B1(n38240), .B2(n36950), .ZN(
        n8019) );
  OAI22_X1 U4539 ( .A1(n38241), .A2(n38687), .B1(n38240), .B2(n36951), .ZN(
        n8020) );
  OAI22_X1 U4540 ( .A1(n38241), .A2(n38694), .B1(n38240), .B2(n36952), .ZN(
        n8021) );
  OAI22_X1 U4541 ( .A1(n38241), .A2(n38701), .B1(n38240), .B2(n36953), .ZN(
        n8022) );
  OAI22_X1 U4542 ( .A1(n38241), .A2(n38708), .B1(n38240), .B2(n36954), .ZN(
        n8023) );
  OAI22_X1 U4543 ( .A1(n38242), .A2(n38715), .B1(n38240), .B2(n36955), .ZN(
        n8024) );
  OAI22_X1 U4544 ( .A1(n38242), .A2(n38722), .B1(n38240), .B2(n36956), .ZN(
        n8025) );
  OAI22_X1 U4545 ( .A1(n38242), .A2(n38729), .B1(n38240), .B2(n36957), .ZN(
        n8026) );
  OAI22_X1 U4546 ( .A1(n38242), .A2(n38736), .B1(n38240), .B2(n36958), .ZN(
        n8027) );
  OAI22_X1 U4547 ( .A1(n38242), .A2(n38743), .B1(n38240), .B2(n36959), .ZN(
        n8028) );
  OAI22_X1 U4548 ( .A1(n38243), .A2(n38750), .B1(n38240), .B2(n36960), .ZN(
        n8029) );
  OAI22_X1 U4549 ( .A1(n38243), .A2(n38757), .B1(n38240), .B2(n36961), .ZN(
        n8030) );
  OAI22_X1 U4550 ( .A1(n38243), .A2(n38764), .B1(n38240), .B2(n36962), .ZN(
        n8031) );
  OAI22_X1 U4551 ( .A1(n38243), .A2(n38771), .B1(n38240), .B2(n36963), .ZN(
        n8032) );
  OAI22_X1 U4552 ( .A1(n38243), .A2(n38778), .B1(n4041), .B2(n36964), .ZN(
        n8033) );
  OAI22_X1 U4553 ( .A1(n38244), .A2(n38785), .B1(n4041), .B2(n36965), .ZN(
        n8034) );
  OAI22_X1 U4554 ( .A1(n38244), .A2(n38792), .B1(n4041), .B2(n36966), .ZN(
        n8035) );
  OAI22_X1 U4555 ( .A1(n38244), .A2(n38799), .B1(n4041), .B2(n36967), .ZN(
        n8036) );
  OAI22_X1 U4556 ( .A1(n38244), .A2(n38806), .B1(n4041), .B2(n36968), .ZN(
        n8037) );
  OAI22_X1 U4557 ( .A1(n38244), .A2(n38813), .B1(n4041), .B2(n36969), .ZN(
        n8038) );
  OAI22_X1 U4558 ( .A1(n38245), .A2(n38820), .B1(n4041), .B2(n36970), .ZN(
        n8039) );
  OAI22_X1 U4559 ( .A1(n38245), .A2(n38827), .B1(n38240), .B2(n36971), .ZN(
        n8040) );
  OAI22_X1 U4560 ( .A1(n38245), .A2(n38834), .B1(n38240), .B2(n36972), .ZN(
        n8041) );
  OAI22_X1 U4561 ( .A1(n38245), .A2(n38841), .B1(n38240), .B2(n36973), .ZN(
        n8042) );
  OAI22_X1 U4562 ( .A1(n38262), .A2(n38680), .B1(n38261), .B2(n37358), .ZN(
        n8083) );
  OAI22_X1 U4563 ( .A1(n38262), .A2(n38687), .B1(n38261), .B2(n37359), .ZN(
        n8084) );
  OAI22_X1 U4564 ( .A1(n38262), .A2(n38694), .B1(n38261), .B2(n37360), .ZN(
        n8085) );
  OAI22_X1 U4565 ( .A1(n38262), .A2(n38701), .B1(n38261), .B2(n37361), .ZN(
        n8086) );
  OAI22_X1 U4566 ( .A1(n38262), .A2(n38708), .B1(n38261), .B2(n37362), .ZN(
        n8087) );
  OAI22_X1 U4567 ( .A1(n38263), .A2(n38715), .B1(n38261), .B2(n37363), .ZN(
        n8088) );
  OAI22_X1 U4568 ( .A1(n38263), .A2(n38722), .B1(n38261), .B2(n37364), .ZN(
        n8089) );
  OAI22_X1 U4569 ( .A1(n38263), .A2(n38729), .B1(n38261), .B2(n37365), .ZN(
        n8090) );
  OAI22_X1 U4570 ( .A1(n38263), .A2(n38736), .B1(n38261), .B2(n37366), .ZN(
        n8091) );
  OAI22_X1 U4571 ( .A1(n38263), .A2(n38743), .B1(n38261), .B2(n37367), .ZN(
        n8092) );
  OAI22_X1 U4572 ( .A1(n38264), .A2(n38750), .B1(n38261), .B2(n37368), .ZN(
        n8093) );
  OAI22_X1 U4573 ( .A1(n38264), .A2(n38757), .B1(n38261), .B2(n37369), .ZN(
        n8094) );
  OAI22_X1 U4574 ( .A1(n38264), .A2(n38764), .B1(n38261), .B2(n37370), .ZN(
        n8095) );
  OAI22_X1 U4575 ( .A1(n38264), .A2(n38771), .B1(n38261), .B2(n37371), .ZN(
        n8096) );
  OAI22_X1 U4576 ( .A1(n38264), .A2(n38778), .B1(n3971), .B2(n37372), .ZN(
        n8097) );
  OAI22_X1 U4577 ( .A1(n38265), .A2(n38785), .B1(n3971), .B2(n37373), .ZN(
        n8098) );
  OAI22_X1 U4578 ( .A1(n38265), .A2(n38792), .B1(n3971), .B2(n37374), .ZN(
        n8099) );
  OAI22_X1 U4579 ( .A1(n38265), .A2(n38799), .B1(n3971), .B2(n37375), .ZN(
        n8100) );
  OAI22_X1 U4580 ( .A1(n38265), .A2(n38806), .B1(n3971), .B2(n37376), .ZN(
        n8101) );
  OAI22_X1 U4581 ( .A1(n38265), .A2(n38813), .B1(n3971), .B2(n37377), .ZN(
        n8102) );
  OAI22_X1 U4582 ( .A1(n38266), .A2(n38820), .B1(n3971), .B2(n37378), .ZN(
        n8103) );
  OAI22_X1 U4583 ( .A1(n38266), .A2(n38827), .B1(n38261), .B2(n37379), .ZN(
        n8104) );
  OAI22_X1 U4584 ( .A1(n38266), .A2(n38834), .B1(n38261), .B2(n37380), .ZN(
        n8105) );
  OAI22_X1 U4585 ( .A1(n38266), .A2(n38841), .B1(n38261), .B2(n37381), .ZN(
        n8106) );
  OAI22_X1 U4586 ( .A1(n38295), .A2(n38680), .B1(n38294), .B2(n36974), .ZN(
        n8179) );
  OAI22_X1 U4587 ( .A1(n38295), .A2(n38687), .B1(n38294), .B2(n36975), .ZN(
        n8180) );
  OAI22_X1 U4588 ( .A1(n38295), .A2(n38694), .B1(n38294), .B2(n36976), .ZN(
        n8181) );
  OAI22_X1 U4589 ( .A1(n38295), .A2(n38701), .B1(n38294), .B2(n36977), .ZN(
        n8182) );
  OAI22_X1 U4590 ( .A1(n38295), .A2(n38708), .B1(n38294), .B2(n36978), .ZN(
        n8183) );
  OAI22_X1 U4591 ( .A1(n38296), .A2(n38715), .B1(n38294), .B2(n36979), .ZN(
        n8184) );
  OAI22_X1 U4592 ( .A1(n38296), .A2(n38722), .B1(n38294), .B2(n36980), .ZN(
        n8185) );
  OAI22_X1 U4593 ( .A1(n38296), .A2(n38729), .B1(n38294), .B2(n36981), .ZN(
        n8186) );
  OAI22_X1 U4594 ( .A1(n38296), .A2(n38736), .B1(n38294), .B2(n36982), .ZN(
        n8187) );
  OAI22_X1 U4595 ( .A1(n38296), .A2(n38743), .B1(n38294), .B2(n36983), .ZN(
        n8188) );
  OAI22_X1 U4596 ( .A1(n38297), .A2(n38750), .B1(n38294), .B2(n36984), .ZN(
        n8189) );
  OAI22_X1 U4597 ( .A1(n38297), .A2(n38757), .B1(n38294), .B2(n36985), .ZN(
        n8190) );
  OAI22_X1 U4598 ( .A1(n38297), .A2(n38764), .B1(n38294), .B2(n36986), .ZN(
        n8191) );
  OAI22_X1 U4599 ( .A1(n38297), .A2(n38771), .B1(n38294), .B2(n36987), .ZN(
        n8192) );
  OAI22_X1 U4600 ( .A1(n38297), .A2(n38778), .B1(n3866), .B2(n36988), .ZN(
        n8193) );
  OAI22_X1 U4601 ( .A1(n38298), .A2(n38785), .B1(n3866), .B2(n36989), .ZN(
        n8194) );
  OAI22_X1 U4602 ( .A1(n38298), .A2(n38792), .B1(n3866), .B2(n36990), .ZN(
        n8195) );
  OAI22_X1 U4603 ( .A1(n38298), .A2(n38799), .B1(n3866), .B2(n36991), .ZN(
        n8196) );
  OAI22_X1 U4604 ( .A1(n38298), .A2(n38806), .B1(n3866), .B2(n36992), .ZN(
        n8197) );
  OAI22_X1 U4605 ( .A1(n38298), .A2(n38813), .B1(n3866), .B2(n36993), .ZN(
        n8198) );
  OAI22_X1 U4606 ( .A1(n38299), .A2(n38820), .B1(n3866), .B2(n36994), .ZN(
        n8199) );
  OAI22_X1 U4607 ( .A1(n38299), .A2(n38827), .B1(n38294), .B2(n36995), .ZN(
        n8200) );
  OAI22_X1 U4608 ( .A1(n38299), .A2(n38834), .B1(n38294), .B2(n36996), .ZN(
        n8201) );
  OAI22_X1 U4609 ( .A1(n38299), .A2(n38841), .B1(n38294), .B2(n36997), .ZN(
        n8202) );
  OAI22_X1 U4610 ( .A1(n38328), .A2(n38679), .B1(n38327), .B2(n36998), .ZN(
        n8275) );
  OAI22_X1 U4611 ( .A1(n38328), .A2(n38686), .B1(n38327), .B2(n36999), .ZN(
        n8276) );
  OAI22_X1 U4612 ( .A1(n38328), .A2(n38693), .B1(n38327), .B2(n37000), .ZN(
        n8277) );
  OAI22_X1 U4613 ( .A1(n38328), .A2(n38700), .B1(n38327), .B2(n37001), .ZN(
        n8278) );
  OAI22_X1 U4614 ( .A1(n38328), .A2(n38707), .B1(n38327), .B2(n37002), .ZN(
        n8279) );
  OAI22_X1 U4615 ( .A1(n38329), .A2(n38714), .B1(n38327), .B2(n37003), .ZN(
        n8280) );
  OAI22_X1 U4616 ( .A1(n38329), .A2(n38721), .B1(n38327), .B2(n37004), .ZN(
        n8281) );
  OAI22_X1 U4617 ( .A1(n38329), .A2(n38728), .B1(n38327), .B2(n37005), .ZN(
        n8282) );
  OAI22_X1 U4618 ( .A1(n38329), .A2(n38735), .B1(n38327), .B2(n37006), .ZN(
        n8283) );
  OAI22_X1 U4619 ( .A1(n38329), .A2(n38742), .B1(n38327), .B2(n37007), .ZN(
        n8284) );
  OAI22_X1 U4620 ( .A1(n38330), .A2(n38749), .B1(n38327), .B2(n37008), .ZN(
        n8285) );
  OAI22_X1 U4621 ( .A1(n38330), .A2(n38756), .B1(n38327), .B2(n37009), .ZN(
        n8286) );
  OAI22_X1 U4622 ( .A1(n38330), .A2(n38763), .B1(n38327), .B2(n37010), .ZN(
        n8287) );
  OAI22_X1 U4623 ( .A1(n38330), .A2(n38770), .B1(n38327), .B2(n37011), .ZN(
        n8288) );
  OAI22_X1 U4624 ( .A1(n38330), .A2(n38777), .B1(n3761), .B2(n37012), .ZN(
        n8289) );
  OAI22_X1 U4625 ( .A1(n38331), .A2(n38784), .B1(n3761), .B2(n37013), .ZN(
        n8290) );
  OAI22_X1 U4626 ( .A1(n38331), .A2(n38791), .B1(n3761), .B2(n37014), .ZN(
        n8291) );
  OAI22_X1 U4627 ( .A1(n38331), .A2(n38798), .B1(n3761), .B2(n37015), .ZN(
        n8292) );
  OAI22_X1 U4628 ( .A1(n38331), .A2(n38805), .B1(n3761), .B2(n37016), .ZN(
        n8293) );
  OAI22_X1 U4629 ( .A1(n38331), .A2(n38812), .B1(n3761), .B2(n37017), .ZN(
        n8294) );
  OAI22_X1 U4630 ( .A1(n38332), .A2(n38819), .B1(n3761), .B2(n37018), .ZN(
        n8295) );
  OAI22_X1 U4631 ( .A1(n38332), .A2(n38826), .B1(n38327), .B2(n37019), .ZN(
        n8296) );
  OAI22_X1 U4632 ( .A1(n38332), .A2(n38833), .B1(n38327), .B2(n37020), .ZN(
        n8297) );
  OAI22_X1 U4633 ( .A1(n38332), .A2(n38840), .B1(n38327), .B2(n37021), .ZN(
        n8298) );
  OAI22_X1 U4634 ( .A1(n38349), .A2(n38679), .B1(n38348), .B2(n37382), .ZN(
        n8339) );
  OAI22_X1 U4635 ( .A1(n38349), .A2(n38686), .B1(n38348), .B2(n37383), .ZN(
        n8340) );
  OAI22_X1 U4636 ( .A1(n38349), .A2(n38693), .B1(n38348), .B2(n37384), .ZN(
        n8341) );
  OAI22_X1 U4637 ( .A1(n38349), .A2(n38700), .B1(n38348), .B2(n37385), .ZN(
        n8342) );
  OAI22_X1 U4638 ( .A1(n38349), .A2(n38707), .B1(n38348), .B2(n37386), .ZN(
        n8343) );
  OAI22_X1 U4639 ( .A1(n38350), .A2(n38714), .B1(n38348), .B2(n37387), .ZN(
        n8344) );
  OAI22_X1 U4640 ( .A1(n38350), .A2(n38721), .B1(n38348), .B2(n37388), .ZN(
        n8345) );
  OAI22_X1 U4641 ( .A1(n38350), .A2(n38728), .B1(n38348), .B2(n37389), .ZN(
        n8346) );
  OAI22_X1 U4642 ( .A1(n38350), .A2(n38735), .B1(n38348), .B2(n37390), .ZN(
        n8347) );
  OAI22_X1 U4643 ( .A1(n38350), .A2(n38742), .B1(n38348), .B2(n37391), .ZN(
        n8348) );
  OAI22_X1 U4644 ( .A1(n38351), .A2(n38749), .B1(n38348), .B2(n37392), .ZN(
        n8349) );
  OAI22_X1 U4645 ( .A1(n38351), .A2(n38756), .B1(n38348), .B2(n37393), .ZN(
        n8350) );
  OAI22_X1 U4646 ( .A1(n38351), .A2(n38763), .B1(n38348), .B2(n37394), .ZN(
        n8351) );
  OAI22_X1 U4647 ( .A1(n38351), .A2(n38770), .B1(n38348), .B2(n37395), .ZN(
        n8352) );
  OAI22_X1 U4648 ( .A1(n38351), .A2(n38777), .B1(n3691), .B2(n37396), .ZN(
        n8353) );
  OAI22_X1 U4649 ( .A1(n38352), .A2(n38784), .B1(n3691), .B2(n37397), .ZN(
        n8354) );
  OAI22_X1 U4650 ( .A1(n38352), .A2(n38791), .B1(n3691), .B2(n37398), .ZN(
        n8355) );
  OAI22_X1 U4651 ( .A1(n38352), .A2(n38798), .B1(n3691), .B2(n37399), .ZN(
        n8356) );
  OAI22_X1 U4652 ( .A1(n38352), .A2(n38805), .B1(n3691), .B2(n37400), .ZN(
        n8357) );
  OAI22_X1 U4653 ( .A1(n38352), .A2(n38812), .B1(n3691), .B2(n37401), .ZN(
        n8358) );
  OAI22_X1 U4654 ( .A1(n38353), .A2(n38819), .B1(n3691), .B2(n37402), .ZN(
        n8359) );
  OAI22_X1 U4655 ( .A1(n38353), .A2(n38826), .B1(n38348), .B2(n37403), .ZN(
        n8360) );
  OAI22_X1 U4656 ( .A1(n38353), .A2(n38833), .B1(n38348), .B2(n37404), .ZN(
        n8361) );
  OAI22_X1 U4657 ( .A1(n38353), .A2(n38840), .B1(n38348), .B2(n37405), .ZN(
        n8362) );
  OAI22_X1 U4658 ( .A1(n38382), .A2(n38679), .B1(n38381), .B2(n37022), .ZN(
        n8435) );
  OAI22_X1 U4659 ( .A1(n38382), .A2(n38686), .B1(n38381), .B2(n37023), .ZN(
        n8436) );
  OAI22_X1 U4660 ( .A1(n38382), .A2(n38693), .B1(n38381), .B2(n37024), .ZN(
        n8437) );
  OAI22_X1 U4661 ( .A1(n38382), .A2(n38700), .B1(n38381), .B2(n37025), .ZN(
        n8438) );
  OAI22_X1 U4662 ( .A1(n38382), .A2(n38707), .B1(n38381), .B2(n37026), .ZN(
        n8439) );
  OAI22_X1 U4663 ( .A1(n38383), .A2(n38714), .B1(n38381), .B2(n37027), .ZN(
        n8440) );
  OAI22_X1 U4664 ( .A1(n38383), .A2(n38721), .B1(n38381), .B2(n37028), .ZN(
        n8441) );
  OAI22_X1 U4665 ( .A1(n38383), .A2(n38728), .B1(n38381), .B2(n37029), .ZN(
        n8442) );
  OAI22_X1 U4666 ( .A1(n38383), .A2(n38735), .B1(n38381), .B2(n37030), .ZN(
        n8443) );
  OAI22_X1 U4667 ( .A1(n38383), .A2(n38742), .B1(n38381), .B2(n37031), .ZN(
        n8444) );
  OAI22_X1 U4668 ( .A1(n38384), .A2(n38749), .B1(n38381), .B2(n37032), .ZN(
        n8445) );
  OAI22_X1 U4669 ( .A1(n38384), .A2(n38756), .B1(n38381), .B2(n37033), .ZN(
        n8446) );
  OAI22_X1 U4670 ( .A1(n38384), .A2(n38763), .B1(n38381), .B2(n37034), .ZN(
        n8447) );
  OAI22_X1 U4671 ( .A1(n38384), .A2(n38770), .B1(n38381), .B2(n37035), .ZN(
        n8448) );
  OAI22_X1 U4672 ( .A1(n38384), .A2(n38777), .B1(n3586), .B2(n37036), .ZN(
        n8449) );
  OAI22_X1 U4673 ( .A1(n38385), .A2(n38784), .B1(n3586), .B2(n37037), .ZN(
        n8450) );
  OAI22_X1 U4674 ( .A1(n38385), .A2(n38791), .B1(n3586), .B2(n37038), .ZN(
        n8451) );
  OAI22_X1 U4675 ( .A1(n38385), .A2(n38798), .B1(n3586), .B2(n37039), .ZN(
        n8452) );
  OAI22_X1 U4676 ( .A1(n38385), .A2(n38805), .B1(n3586), .B2(n37040), .ZN(
        n8453) );
  OAI22_X1 U4677 ( .A1(n38385), .A2(n38812), .B1(n3586), .B2(n37041), .ZN(
        n8454) );
  OAI22_X1 U4678 ( .A1(n38386), .A2(n38819), .B1(n3586), .B2(n37042), .ZN(
        n8455) );
  OAI22_X1 U4679 ( .A1(n38386), .A2(n38826), .B1(n38381), .B2(n37043), .ZN(
        n8456) );
  OAI22_X1 U4680 ( .A1(n38386), .A2(n38833), .B1(n38381), .B2(n37044), .ZN(
        n8457) );
  OAI22_X1 U4681 ( .A1(n38386), .A2(n38840), .B1(n38381), .B2(n37045), .ZN(
        n8458) );
  OAI22_X1 U4682 ( .A1(n38403), .A2(n38679), .B1(n38402), .B2(n37406), .ZN(
        n8499) );
  OAI22_X1 U4683 ( .A1(n38403), .A2(n38686), .B1(n38402), .B2(n37407), .ZN(
        n8500) );
  OAI22_X1 U4684 ( .A1(n38403), .A2(n38693), .B1(n38402), .B2(n37408), .ZN(
        n8501) );
  OAI22_X1 U4685 ( .A1(n38403), .A2(n38700), .B1(n38402), .B2(n37409), .ZN(
        n8502) );
  OAI22_X1 U4686 ( .A1(n38403), .A2(n38707), .B1(n38402), .B2(n37410), .ZN(
        n8503) );
  OAI22_X1 U4687 ( .A1(n38404), .A2(n38714), .B1(n38402), .B2(n37411), .ZN(
        n8504) );
  OAI22_X1 U4688 ( .A1(n38404), .A2(n38721), .B1(n38402), .B2(n37412), .ZN(
        n8505) );
  OAI22_X1 U4689 ( .A1(n38404), .A2(n38728), .B1(n38402), .B2(n37413), .ZN(
        n8506) );
  OAI22_X1 U4690 ( .A1(n38404), .A2(n38735), .B1(n38402), .B2(n37414), .ZN(
        n8507) );
  OAI22_X1 U4691 ( .A1(n38404), .A2(n38742), .B1(n38402), .B2(n37415), .ZN(
        n8508) );
  OAI22_X1 U4692 ( .A1(n38405), .A2(n38749), .B1(n38402), .B2(n37416), .ZN(
        n8509) );
  OAI22_X1 U4693 ( .A1(n38405), .A2(n38756), .B1(n38402), .B2(n37417), .ZN(
        n8510) );
  OAI22_X1 U4694 ( .A1(n38405), .A2(n38763), .B1(n38402), .B2(n37418), .ZN(
        n8511) );
  OAI22_X1 U4695 ( .A1(n38405), .A2(n38770), .B1(n38402), .B2(n37419), .ZN(
        n8512) );
  OAI22_X1 U4696 ( .A1(n38405), .A2(n38777), .B1(n3516), .B2(n37420), .ZN(
        n8513) );
  OAI22_X1 U4697 ( .A1(n38406), .A2(n38784), .B1(n3516), .B2(n37421), .ZN(
        n8514) );
  OAI22_X1 U4698 ( .A1(n38406), .A2(n38791), .B1(n3516), .B2(n37422), .ZN(
        n8515) );
  OAI22_X1 U4699 ( .A1(n38406), .A2(n38798), .B1(n3516), .B2(n37423), .ZN(
        n8516) );
  OAI22_X1 U4700 ( .A1(n38406), .A2(n38805), .B1(n3516), .B2(n37424), .ZN(
        n8517) );
  OAI22_X1 U4701 ( .A1(n38406), .A2(n38812), .B1(n3516), .B2(n37425), .ZN(
        n8518) );
  OAI22_X1 U4702 ( .A1(n38407), .A2(n38819), .B1(n3516), .B2(n37426), .ZN(
        n8519) );
  OAI22_X1 U4703 ( .A1(n38407), .A2(n38826), .B1(n38402), .B2(n37427), .ZN(
        n8520) );
  OAI22_X1 U4704 ( .A1(n38407), .A2(n38833), .B1(n38402), .B2(n37428), .ZN(
        n8521) );
  OAI22_X1 U4705 ( .A1(n38407), .A2(n38840), .B1(n38402), .B2(n37429), .ZN(
        n8522) );
  OAI22_X1 U4706 ( .A1(n38436), .A2(n38679), .B1(n38435), .B2(n37046), .ZN(
        n8595) );
  OAI22_X1 U4707 ( .A1(n38436), .A2(n38686), .B1(n38435), .B2(n37047), .ZN(
        n8596) );
  OAI22_X1 U4708 ( .A1(n38436), .A2(n38693), .B1(n38435), .B2(n37048), .ZN(
        n8597) );
  OAI22_X1 U4709 ( .A1(n38436), .A2(n38700), .B1(n38435), .B2(n37049), .ZN(
        n8598) );
  OAI22_X1 U4710 ( .A1(n38436), .A2(n38707), .B1(n38435), .B2(n37050), .ZN(
        n8599) );
  OAI22_X1 U4711 ( .A1(n38437), .A2(n38714), .B1(n38435), .B2(n37051), .ZN(
        n8600) );
  OAI22_X1 U4712 ( .A1(n38437), .A2(n38721), .B1(n38435), .B2(n37052), .ZN(
        n8601) );
  OAI22_X1 U4713 ( .A1(n38437), .A2(n38728), .B1(n38435), .B2(n37053), .ZN(
        n8602) );
  OAI22_X1 U4714 ( .A1(n38437), .A2(n38735), .B1(n38435), .B2(n37054), .ZN(
        n8603) );
  OAI22_X1 U4715 ( .A1(n38437), .A2(n38742), .B1(n38435), .B2(n37055), .ZN(
        n8604) );
  OAI22_X1 U4716 ( .A1(n38438), .A2(n38749), .B1(n38435), .B2(n37056), .ZN(
        n8605) );
  OAI22_X1 U4717 ( .A1(n38438), .A2(n38756), .B1(n38435), .B2(n37057), .ZN(
        n8606) );
  OAI22_X1 U4718 ( .A1(n38438), .A2(n38763), .B1(n38435), .B2(n37058), .ZN(
        n8607) );
  OAI22_X1 U4719 ( .A1(n38438), .A2(n38770), .B1(n38435), .B2(n37059), .ZN(
        n8608) );
  OAI22_X1 U4720 ( .A1(n38438), .A2(n38777), .B1(n3411), .B2(n37060), .ZN(
        n8609) );
  OAI22_X1 U4721 ( .A1(n38439), .A2(n38784), .B1(n3411), .B2(n37061), .ZN(
        n8610) );
  OAI22_X1 U4722 ( .A1(n38439), .A2(n38791), .B1(n3411), .B2(n37062), .ZN(
        n8611) );
  OAI22_X1 U4723 ( .A1(n38439), .A2(n38798), .B1(n3411), .B2(n37063), .ZN(
        n8612) );
  OAI22_X1 U4724 ( .A1(n38439), .A2(n38805), .B1(n3411), .B2(n37064), .ZN(
        n8613) );
  OAI22_X1 U4725 ( .A1(n38439), .A2(n38812), .B1(n3411), .B2(n37065), .ZN(
        n8614) );
  OAI22_X1 U4726 ( .A1(n38440), .A2(n38819), .B1(n3411), .B2(n37066), .ZN(
        n8615) );
  OAI22_X1 U4727 ( .A1(n38440), .A2(n38826), .B1(n38435), .B2(n37067), .ZN(
        n8616) );
  OAI22_X1 U4728 ( .A1(n38440), .A2(n38833), .B1(n38435), .B2(n37068), .ZN(
        n8617) );
  OAI22_X1 U4729 ( .A1(n38440), .A2(n38840), .B1(n38435), .B2(n37069), .ZN(
        n8618) );
  OAI22_X1 U4730 ( .A1(n38457), .A2(n38678), .B1(n38456), .B2(n37430), .ZN(
        n8659) );
  OAI22_X1 U4731 ( .A1(n38457), .A2(n38685), .B1(n38456), .B2(n37431), .ZN(
        n8660) );
  OAI22_X1 U4732 ( .A1(n38457), .A2(n38692), .B1(n38456), .B2(n37432), .ZN(
        n8661) );
  OAI22_X1 U4733 ( .A1(n38457), .A2(n38699), .B1(n38456), .B2(n37433), .ZN(
        n8662) );
  OAI22_X1 U4734 ( .A1(n38457), .A2(n38706), .B1(n38456), .B2(n37434), .ZN(
        n8663) );
  OAI22_X1 U4735 ( .A1(n38458), .A2(n38713), .B1(n38456), .B2(n37435), .ZN(
        n8664) );
  OAI22_X1 U4736 ( .A1(n38458), .A2(n38720), .B1(n38456), .B2(n37436), .ZN(
        n8665) );
  OAI22_X1 U4737 ( .A1(n38458), .A2(n38727), .B1(n38456), .B2(n37437), .ZN(
        n8666) );
  OAI22_X1 U4738 ( .A1(n38458), .A2(n38734), .B1(n38456), .B2(n37438), .ZN(
        n8667) );
  OAI22_X1 U4739 ( .A1(n38458), .A2(n38741), .B1(n38456), .B2(n37439), .ZN(
        n8668) );
  OAI22_X1 U4740 ( .A1(n38459), .A2(n38748), .B1(n38456), .B2(n37440), .ZN(
        n8669) );
  OAI22_X1 U4741 ( .A1(n38459), .A2(n38755), .B1(n38456), .B2(n37441), .ZN(
        n8670) );
  OAI22_X1 U4742 ( .A1(n38459), .A2(n38762), .B1(n38456), .B2(n37442), .ZN(
        n8671) );
  OAI22_X1 U4743 ( .A1(n38459), .A2(n38769), .B1(n38456), .B2(n37443), .ZN(
        n8672) );
  OAI22_X1 U4744 ( .A1(n38459), .A2(n38776), .B1(n3341), .B2(n37444), .ZN(
        n8673) );
  OAI22_X1 U4745 ( .A1(n38460), .A2(n38783), .B1(n3341), .B2(n37445), .ZN(
        n8674) );
  OAI22_X1 U4746 ( .A1(n38460), .A2(n38790), .B1(n3341), .B2(n37446), .ZN(
        n8675) );
  OAI22_X1 U4747 ( .A1(n38460), .A2(n38797), .B1(n3341), .B2(n37447), .ZN(
        n8676) );
  OAI22_X1 U4748 ( .A1(n38460), .A2(n38804), .B1(n3341), .B2(n37448), .ZN(
        n8677) );
  OAI22_X1 U4749 ( .A1(n38460), .A2(n38811), .B1(n3341), .B2(n37449), .ZN(
        n8678) );
  OAI22_X1 U4750 ( .A1(n38461), .A2(n38818), .B1(n3341), .B2(n37450), .ZN(
        n8679) );
  OAI22_X1 U4751 ( .A1(n38461), .A2(n38825), .B1(n38456), .B2(n37451), .ZN(
        n8680) );
  OAI22_X1 U4752 ( .A1(n38461), .A2(n38832), .B1(n38456), .B2(n37452), .ZN(
        n8681) );
  OAI22_X1 U4753 ( .A1(n38461), .A2(n38839), .B1(n38456), .B2(n37453), .ZN(
        n8682) );
  OAI22_X1 U4754 ( .A1(n4083), .A2(n37785), .B1(n9561), .B2(n37794), .ZN(n6675) );
  NOR4_X1 U4755 ( .A1(n9562), .A2(n9563), .A3(n9564), .A4(n9565), .ZN(n9561)
         );
  NAND4_X1 U4756 ( .A1(n9620), .A2(n9621), .A3(n9622), .A4(n9623), .ZN(n9562)
         );
  NAND4_X1 U4757 ( .A1(n9607), .A2(n9608), .A3(n9610), .A4(n9611), .ZN(n9563)
         );
  OAI22_X1 U4758 ( .A1(n4085), .A2(n37785), .B1(n9518), .B2(n37794), .ZN(n6677) );
  NOR4_X1 U4759 ( .A1(n9519), .A2(n9520), .A3(n9521), .A4(n9522), .ZN(n9518)
         );
  NAND4_X1 U4760 ( .A1(n9551), .A2(n9552), .A3(n9553), .A4(n9554), .ZN(n9519)
         );
  NAND4_X1 U4761 ( .A1(n9539), .A2(n9540), .A3(n9541), .A4(n9543), .ZN(n9520)
         );
  OAI22_X1 U4762 ( .A1(n4087), .A2(n37785), .B1(n9476), .B2(n37794), .ZN(n6679) );
  NOR4_X1 U4763 ( .A1(n9477), .A2(n9478), .A3(n9479), .A4(n9480), .ZN(n9476)
         );
  NAND4_X1 U4764 ( .A1(n9509), .A2(n9510), .A3(n9511), .A4(n9512), .ZN(n9477)
         );
  NAND4_X1 U4765 ( .A1(n9497), .A2(n9498), .A3(n9499), .A4(n9501), .ZN(n9478)
         );
  OAI22_X1 U4766 ( .A1(n4089), .A2(n37785), .B1(n9434), .B2(n37794), .ZN(n6681) );
  NOR4_X1 U4767 ( .A1(n9435), .A2(n9436), .A3(n9437), .A4(n9438), .ZN(n9434)
         );
  NAND4_X1 U4768 ( .A1(n9467), .A2(n9468), .A3(n9469), .A4(n9470), .ZN(n9435)
         );
  NAND4_X1 U4769 ( .A1(n9455), .A2(n9456), .A3(n9457), .A4(n9459), .ZN(n9436)
         );
  OAI22_X1 U4770 ( .A1(n4091), .A2(n37785), .B1(n9392), .B2(n37793), .ZN(n6683) );
  NOR4_X1 U4771 ( .A1(n9393), .A2(n9394), .A3(n9395), .A4(n9396), .ZN(n9392)
         );
  NAND4_X1 U4772 ( .A1(n9425), .A2(n9426), .A3(n9427), .A4(n9428), .ZN(n9393)
         );
  NAND4_X1 U4773 ( .A1(n9413), .A2(n9414), .A3(n9415), .A4(n9417), .ZN(n9394)
         );
  OAI22_X1 U4774 ( .A1(n4093), .A2(n37785), .B1(n9350), .B2(n37793), .ZN(n6685) );
  NOR4_X1 U4775 ( .A1(n9351), .A2(n9352), .A3(n9353), .A4(n9354), .ZN(n9350)
         );
  NAND4_X1 U4776 ( .A1(n9383), .A2(n9384), .A3(n9385), .A4(n9386), .ZN(n9351)
         );
  NAND4_X1 U4777 ( .A1(n9371), .A2(n9372), .A3(n9373), .A4(n9375), .ZN(n9352)
         );
  OAI22_X1 U4778 ( .A1(n4095), .A2(n37785), .B1(n9308), .B2(n37793), .ZN(n6687) );
  NOR4_X1 U4779 ( .A1(n9309), .A2(n9310), .A3(n9311), .A4(n9312), .ZN(n9308)
         );
  NAND4_X1 U4780 ( .A1(n9341), .A2(n9342), .A3(n9343), .A4(n9344), .ZN(n9309)
         );
  NAND4_X1 U4781 ( .A1(n9329), .A2(n9330), .A3(n9331), .A4(n9333), .ZN(n9310)
         );
  OAI22_X1 U4782 ( .A1(n4097), .A2(n37785), .B1(n6674), .B2(n37793), .ZN(n6689) );
  NOR4_X1 U4783 ( .A1(n9267), .A2(n9268), .A3(n9269), .A4(n9270), .ZN(n6674)
         );
  NAND4_X1 U4784 ( .A1(n9299), .A2(n9300), .A3(n9301), .A4(n9302), .ZN(n9267)
         );
  NAND4_X1 U4785 ( .A1(n9287), .A2(n9288), .A3(n9289), .A4(n9291), .ZN(n9268)
         );
  OAI22_X1 U4786 ( .A1(n4099), .A2(n37785), .B1(n6632), .B2(n37792), .ZN(n6691) );
  NOR4_X1 U4787 ( .A1(n6633), .A2(n6634), .A3(n6635), .A4(n6636), .ZN(n6632)
         );
  NAND4_X1 U4788 ( .A1(n6665), .A2(n6666), .A3(n6667), .A4(n6668), .ZN(n6633)
         );
  NAND4_X1 U4789 ( .A1(n6653), .A2(n6654), .A3(n6655), .A4(n6657), .ZN(n6634)
         );
  OAI22_X1 U4790 ( .A1(n4101), .A2(n37785), .B1(n6590), .B2(n37792), .ZN(n6693) );
  NOR4_X1 U4791 ( .A1(n6591), .A2(n6592), .A3(n6593), .A4(n6594), .ZN(n6590)
         );
  NAND4_X1 U4792 ( .A1(n6623), .A2(n6624), .A3(n6625), .A4(n6626), .ZN(n6591)
         );
  NAND4_X1 U4793 ( .A1(n6611), .A2(n6612), .A3(n6613), .A4(n6615), .ZN(n6592)
         );
  OAI22_X1 U4794 ( .A1(n4103), .A2(n37785), .B1(n6548), .B2(n37792), .ZN(n6695) );
  NOR4_X1 U4795 ( .A1(n6549), .A2(n6550), .A3(n6551), .A4(n6552), .ZN(n6548)
         );
  NAND4_X1 U4796 ( .A1(n6581), .A2(n6582), .A3(n6583), .A4(n6584), .ZN(n6549)
         );
  NAND4_X1 U4797 ( .A1(n6569), .A2(n6570), .A3(n6571), .A4(n6573), .ZN(n6550)
         );
  OAI22_X1 U4798 ( .A1(n4105), .A2(n37785), .B1(n6482), .B2(n37792), .ZN(n6697) );
  NOR4_X1 U4799 ( .A1(n6484), .A2(n6508), .A3(n6509), .A4(n6510), .ZN(n6482)
         );
  NAND4_X1 U4800 ( .A1(n6539), .A2(n6540), .A3(n6541), .A4(n6542), .ZN(n6484)
         );
  NAND4_X1 U4801 ( .A1(n6527), .A2(n6528), .A3(n6529), .A4(n6531), .ZN(n6508)
         );
  OAI22_X1 U4802 ( .A1(n4107), .A2(n37786), .B1(n6336), .B2(n37791), .ZN(n6699) );
  NOR4_X1 U4803 ( .A1(n6337), .A2(n6338), .A3(n6339), .A4(n6340), .ZN(n6336)
         );
  NAND4_X1 U4804 ( .A1(n6373), .A2(n6406), .A3(n6408), .A4(n6441), .ZN(n6337)
         );
  NAND4_X1 U4805 ( .A1(n6357), .A2(n6358), .A3(n6359), .A4(n6361), .ZN(n6338)
         );
  OAI22_X1 U4806 ( .A1(n4109), .A2(n37786), .B1(n6294), .B2(n37791), .ZN(n6701) );
  NOR4_X1 U4807 ( .A1(n6295), .A2(n6296), .A3(n6297), .A4(n6298), .ZN(n6294)
         );
  NAND4_X1 U4808 ( .A1(n6327), .A2(n6328), .A3(n6329), .A4(n6330), .ZN(n6295)
         );
  NAND4_X1 U4809 ( .A1(n6315), .A2(n6316), .A3(n6317), .A4(n6319), .ZN(n6296)
         );
  OAI22_X1 U4810 ( .A1(n4111), .A2(n37786), .B1(n6252), .B2(n37791), .ZN(n6703) );
  NOR4_X1 U4811 ( .A1(n6253), .A2(n6254), .A3(n6255), .A4(n6256), .ZN(n6252)
         );
  NAND4_X1 U4812 ( .A1(n6285), .A2(n6286), .A3(n6287), .A4(n6288), .ZN(n6253)
         );
  NAND4_X1 U4813 ( .A1(n6273), .A2(n6274), .A3(n6275), .A4(n6277), .ZN(n6254)
         );
  OAI22_X1 U4814 ( .A1(n4113), .A2(n37786), .B1(n6210), .B2(n37791), .ZN(n6705) );
  NOR4_X1 U4815 ( .A1(n6211), .A2(n6212), .A3(n6213), .A4(n6214), .ZN(n6210)
         );
  NAND4_X1 U4816 ( .A1(n6243), .A2(n6244), .A3(n6245), .A4(n6246), .ZN(n6211)
         );
  NAND4_X1 U4817 ( .A1(n6231), .A2(n6232), .A3(n6233), .A4(n6235), .ZN(n6212)
         );
  OAI22_X1 U4818 ( .A1(n4115), .A2(n37786), .B1(n6168), .B2(n37790), .ZN(n6707) );
  NOR4_X1 U4819 ( .A1(n6169), .A2(n6170), .A3(n6171), .A4(n6172), .ZN(n6168)
         );
  NAND4_X1 U4820 ( .A1(n6201), .A2(n6202), .A3(n6203), .A4(n6204), .ZN(n6169)
         );
  NAND4_X1 U4821 ( .A1(n6189), .A2(n6190), .A3(n6191), .A4(n6193), .ZN(n6170)
         );
  OAI22_X1 U4822 ( .A1(n4117), .A2(n37786), .B1(n6126), .B2(n37790), .ZN(n6709) );
  NOR4_X1 U4823 ( .A1(n6127), .A2(n6128), .A3(n6129), .A4(n6130), .ZN(n6126)
         );
  NAND4_X1 U4824 ( .A1(n6159), .A2(n6160), .A3(n6161), .A4(n6162), .ZN(n6127)
         );
  NAND4_X1 U4825 ( .A1(n6147), .A2(n6148), .A3(n6149), .A4(n6151), .ZN(n6128)
         );
  OAI22_X1 U4826 ( .A1(n4119), .A2(n37786), .B1(n6084), .B2(n37790), .ZN(n6711) );
  NOR4_X1 U4827 ( .A1(n6085), .A2(n6086), .A3(n6087), .A4(n6088), .ZN(n6084)
         );
  NAND4_X1 U4828 ( .A1(n6117), .A2(n6118), .A3(n6119), .A4(n6120), .ZN(n6085)
         );
  NAND4_X1 U4829 ( .A1(n6105), .A2(n6106), .A3(n6107), .A4(n6109), .ZN(n6086)
         );
  OAI22_X1 U4830 ( .A1(n4121), .A2(n37786), .B1(n6042), .B2(n37790), .ZN(n6713) );
  NOR4_X1 U4831 ( .A1(n6043), .A2(n6044), .A3(n6045), .A4(n6046), .ZN(n6042)
         );
  NAND4_X1 U4832 ( .A1(n6075), .A2(n6076), .A3(n6077), .A4(n6078), .ZN(n6043)
         );
  NAND4_X1 U4833 ( .A1(n6063), .A2(n6064), .A3(n6065), .A4(n6067), .ZN(n6044)
         );
  OAI22_X1 U4834 ( .A1(n4123), .A2(n37786), .B1(n6000), .B2(n37789), .ZN(n6715) );
  NOR4_X1 U4835 ( .A1(n6001), .A2(n6002), .A3(n6003), .A4(n6004), .ZN(n6000)
         );
  NAND4_X1 U4836 ( .A1(n6033), .A2(n6034), .A3(n6035), .A4(n6036), .ZN(n6001)
         );
  NAND4_X1 U4837 ( .A1(n6021), .A2(n6022), .A3(n6023), .A4(n6025), .ZN(n6002)
         );
  OAI22_X1 U4838 ( .A1(n4125), .A2(n37786), .B1(n5958), .B2(n37789), .ZN(n6717) );
  NOR4_X1 U4839 ( .A1(n5959), .A2(n5960), .A3(n5961), .A4(n5962), .ZN(n5958)
         );
  NAND4_X1 U4840 ( .A1(n5991), .A2(n5992), .A3(n5993), .A4(n5994), .ZN(n5959)
         );
  NAND4_X1 U4841 ( .A1(n5979), .A2(n5980), .A3(n5981), .A4(n5983), .ZN(n5960)
         );
  OAI22_X1 U4842 ( .A1(n4127), .A2(n37786), .B1(n5916), .B2(n37789), .ZN(n6719) );
  NOR4_X1 U4843 ( .A1(n5917), .A2(n5918), .A3(n5919), .A4(n5920), .ZN(n5916)
         );
  NAND4_X1 U4844 ( .A1(n5949), .A2(n5950), .A3(n5951), .A4(n5952), .ZN(n5917)
         );
  NAND4_X1 U4845 ( .A1(n5937), .A2(n5938), .A3(n5939), .A4(n5941), .ZN(n5918)
         );
  OAI22_X1 U4846 ( .A1(n4129), .A2(n37786), .B1(n5874), .B2(n37789), .ZN(n6721) );
  NOR4_X1 U4847 ( .A1(n5875), .A2(n5876), .A3(n5877), .A4(n5878), .ZN(n5874)
         );
  NAND4_X1 U4848 ( .A1(n5907), .A2(n5908), .A3(n5909), .A4(n5910), .ZN(n5875)
         );
  NAND4_X1 U4849 ( .A1(n5895), .A2(n5896), .A3(n5897), .A4(n5899), .ZN(n5876)
         );
  OAI22_X1 U4850 ( .A1(n4131), .A2(n37785), .B1(n5832), .B2(n37788), .ZN(n6723) );
  NOR4_X1 U4851 ( .A1(n5833), .A2(n5834), .A3(n5835), .A4(n5836), .ZN(n5832)
         );
  NAND4_X1 U4852 ( .A1(n5865), .A2(n5866), .A3(n5867), .A4(n5868), .ZN(n5833)
         );
  NAND4_X1 U4853 ( .A1(n5853), .A2(n5854), .A3(n5855), .A4(n5857), .ZN(n5834)
         );
  OAI22_X1 U4854 ( .A1(n4133), .A2(n37786), .B1(n5790), .B2(n37788), .ZN(n6725) );
  NOR4_X1 U4855 ( .A1(n5791), .A2(n5792), .A3(n5793), .A4(n5794), .ZN(n5790)
         );
  NAND4_X1 U4856 ( .A1(n5823), .A2(n5824), .A3(n5825), .A4(n5826), .ZN(n5791)
         );
  NAND4_X1 U4857 ( .A1(n5811), .A2(n5812), .A3(n5813), .A4(n5815), .ZN(n5792)
         );
  OAI22_X1 U4858 ( .A1(n4135), .A2(n37785), .B1(n5748), .B2(n37788), .ZN(n6727) );
  NOR4_X1 U4859 ( .A1(n5749), .A2(n5750), .A3(n5751), .A4(n5752), .ZN(n5748)
         );
  NAND4_X1 U4860 ( .A1(n5781), .A2(n5782), .A3(n5783), .A4(n5784), .ZN(n5749)
         );
  NAND4_X1 U4861 ( .A1(n5769), .A2(n5770), .A3(n5771), .A4(n5773), .ZN(n5750)
         );
  OAI22_X1 U4862 ( .A1(n4137), .A2(n37786), .B1(n5706), .B2(n37788), .ZN(n6729) );
  NOR4_X1 U4863 ( .A1(n5707), .A2(n5708), .A3(n5709), .A4(n5710), .ZN(n5706)
         );
  NAND4_X1 U4864 ( .A1(n5739), .A2(n5740), .A3(n5741), .A4(n5742), .ZN(n5707)
         );
  NAND4_X1 U4865 ( .A1(n5727), .A2(n5728), .A3(n5729), .A4(n5731), .ZN(n5708)
         );
  OAI22_X1 U4866 ( .A1(n4139), .A2(n37785), .B1(n5664), .B2(n37787), .ZN(n6731) );
  NOR4_X1 U4867 ( .A1(n5665), .A2(n5666), .A3(n5667), .A4(n5668), .ZN(n5664)
         );
  NAND4_X1 U4868 ( .A1(n5697), .A2(n5698), .A3(n5699), .A4(n5700), .ZN(n5665)
         );
  NAND4_X1 U4869 ( .A1(n5685), .A2(n5686), .A3(n5687), .A4(n5689), .ZN(n5666)
         );
  OAI22_X1 U4870 ( .A1(n4141), .A2(n37786), .B1(n5622), .B2(n37787), .ZN(n6733) );
  NOR4_X1 U4871 ( .A1(n5623), .A2(n5624), .A3(n5625), .A4(n5626), .ZN(n5622)
         );
  NAND4_X1 U4872 ( .A1(n5655), .A2(n5656), .A3(n5657), .A4(n5658), .ZN(n5623)
         );
  NAND4_X1 U4873 ( .A1(n5643), .A2(n5644), .A3(n5645), .A4(n5647), .ZN(n5624)
         );
  OAI22_X1 U4874 ( .A1(n4143), .A2(n37785), .B1(n5580), .B2(n37787), .ZN(n6735) );
  NOR4_X1 U4875 ( .A1(n5581), .A2(n5582), .A3(n5583), .A4(n5584), .ZN(n5580)
         );
  NAND4_X1 U4876 ( .A1(n5613), .A2(n5614), .A3(n5615), .A4(n5616), .ZN(n5581)
         );
  NAND4_X1 U4877 ( .A1(n5601), .A2(n5602), .A3(n5603), .A4(n5605), .ZN(n5582)
         );
  OAI22_X1 U4878 ( .A1(n4145), .A2(n37786), .B1(n5512), .B2(n37787), .ZN(n6737) );
  NOR4_X1 U4879 ( .A1(n5514), .A2(n5515), .A3(n5516), .A4(n5517), .ZN(n5512)
         );
  NAND4_X1 U4880 ( .A1(n5563), .A2(n5564), .A3(n5565), .A4(n5566), .ZN(n5514)
         );
  NAND4_X1 U4881 ( .A1(n5543), .A2(n5544), .A3(n5545), .A4(n5546), .ZN(n5515)
         );
  NAND4_X1 U4882 ( .A1(n9566), .A2(n9567), .A3(n9568), .A4(n9569), .ZN(n9565)
         );
  AOI221_X1 U4883 ( .B1(net253583), .B2(n37764), .C1(net253551), .C2(n37761), 
        .A(n9588), .ZN(n9566) );
  AOI221_X1 U4884 ( .B1(net253903), .B2(n37770), .C1(net254095), .C2(n37767), 
        .A(n9582), .ZN(n9567) );
  AOI221_X1 U4885 ( .B1(net253711), .B2(n37776), .C1(net253679), .C2(n37773), 
        .A(n9576), .ZN(n9568) );
  NAND4_X1 U4886 ( .A1(n9523), .A2(n9524), .A3(n9525), .A4(n9526), .ZN(n9522)
         );
  AOI221_X1 U4887 ( .B1(net253584), .B2(n37764), .C1(net253552), .C2(n37761), 
        .A(n9530), .ZN(n9523) );
  AOI221_X1 U4888 ( .B1(net253904), .B2(n37770), .C1(net254096), .C2(n37767), 
        .A(n9529), .ZN(n9524) );
  AOI221_X1 U4889 ( .B1(net253712), .B2(n37776), .C1(net253680), .C2(n37773), 
        .A(n9528), .ZN(n9525) );
  NAND4_X1 U4890 ( .A1(n9481), .A2(n9482), .A3(n9483), .A4(n9484), .ZN(n9480)
         );
  AOI221_X1 U4891 ( .B1(net253585), .B2(n37764), .C1(net253553), .C2(n37761), 
        .A(n9488), .ZN(n9481) );
  AOI221_X1 U4892 ( .B1(net253905), .B2(n37770), .C1(net254097), .C2(n37767), 
        .A(n9487), .ZN(n9482) );
  AOI221_X1 U4893 ( .B1(net253713), .B2(n37776), .C1(net253681), .C2(n37773), 
        .A(n9486), .ZN(n9483) );
  NAND4_X1 U4894 ( .A1(n9439), .A2(n9440), .A3(n9441), .A4(n9442), .ZN(n9438)
         );
  AOI221_X1 U4895 ( .B1(net253586), .B2(n37764), .C1(net253554), .C2(n37761), 
        .A(n9446), .ZN(n9439) );
  AOI221_X1 U4896 ( .B1(net253906), .B2(n37770), .C1(net254098), .C2(n37767), 
        .A(n9445), .ZN(n9440) );
  AOI221_X1 U4897 ( .B1(net253714), .B2(n37776), .C1(net253682), .C2(n37773), 
        .A(n9444), .ZN(n9441) );
  NAND4_X1 U4898 ( .A1(n9397), .A2(n9398), .A3(n9399), .A4(n9400), .ZN(n9396)
         );
  AOI221_X1 U4899 ( .B1(net253587), .B2(n37764), .C1(net253555), .C2(n37761), 
        .A(n9404), .ZN(n9397) );
  AOI221_X1 U4900 ( .B1(net253907), .B2(n37770), .C1(net254099), .C2(n37767), 
        .A(n9403), .ZN(n9398) );
  AOI221_X1 U4901 ( .B1(net253715), .B2(n37776), .C1(net253683), .C2(n37773), 
        .A(n9402), .ZN(n9399) );
  NAND4_X1 U4902 ( .A1(n9355), .A2(n9356), .A3(n9357), .A4(n9358), .ZN(n9354)
         );
  AOI221_X1 U4903 ( .B1(net253588), .B2(n37764), .C1(net253556), .C2(n37761), 
        .A(n9362), .ZN(n9355) );
  AOI221_X1 U4904 ( .B1(net253908), .B2(n37770), .C1(net254100), .C2(n37767), 
        .A(n9361), .ZN(n9356) );
  AOI221_X1 U4905 ( .B1(net253716), .B2(n37776), .C1(net253684), .C2(n37773), 
        .A(n9360), .ZN(n9357) );
  NAND4_X1 U4906 ( .A1(n9313), .A2(n9314), .A3(n9315), .A4(n9316), .ZN(n9312)
         );
  AOI221_X1 U4907 ( .B1(net253589), .B2(n37764), .C1(net253557), .C2(n37761), 
        .A(n9320), .ZN(n9313) );
  AOI221_X1 U4908 ( .B1(net253909), .B2(n37770), .C1(net254101), .C2(n37767), 
        .A(n9319), .ZN(n9314) );
  AOI221_X1 U4909 ( .B1(net253717), .B2(n37776), .C1(net253685), .C2(n37773), 
        .A(n9318), .ZN(n9315) );
  NAND4_X1 U4910 ( .A1(n9271), .A2(n9272), .A3(n9273), .A4(n9274), .ZN(n9270)
         );
  AOI221_X1 U4911 ( .B1(net253590), .B2(n37764), .C1(net253558), .C2(n37761), 
        .A(n9278), .ZN(n9271) );
  AOI221_X1 U4912 ( .B1(net253910), .B2(n37770), .C1(net254102), .C2(n37767), 
        .A(n9277), .ZN(n9272) );
  AOI221_X1 U4913 ( .B1(net253718), .B2(n37776), .C1(net253686), .C2(n37773), 
        .A(n9276), .ZN(n9273) );
  NAND4_X1 U4914 ( .A1(n6637), .A2(n6638), .A3(n6639), .A4(n6640), .ZN(n6636)
         );
  AOI221_X1 U4915 ( .B1(net253591), .B2(n37764), .C1(net253559), .C2(n37761), 
        .A(n6644), .ZN(n6637) );
  AOI221_X1 U4916 ( .B1(net253911), .B2(n37770), .C1(net254103), .C2(n37767), 
        .A(n6643), .ZN(n6638) );
  AOI221_X1 U4917 ( .B1(net253719), .B2(n37776), .C1(net253687), .C2(n37773), 
        .A(n6642), .ZN(n6639) );
  NAND4_X1 U4918 ( .A1(n6595), .A2(n6596), .A3(n6597), .A4(n6598), .ZN(n6594)
         );
  AOI221_X1 U4919 ( .B1(net253592), .B2(n37764), .C1(net253560), .C2(n37761), 
        .A(n6602), .ZN(n6595) );
  AOI221_X1 U4920 ( .B1(net253912), .B2(n37770), .C1(net254104), .C2(n37767), 
        .A(n6601), .ZN(n6596) );
  AOI221_X1 U4921 ( .B1(net253720), .B2(n37776), .C1(net253688), .C2(n37773), 
        .A(n6600), .ZN(n6597) );
  NAND4_X1 U4922 ( .A1(n6553), .A2(n6554), .A3(n6555), .A4(n6556), .ZN(n6552)
         );
  AOI221_X1 U4923 ( .B1(net253593), .B2(n37764), .C1(net253561), .C2(n37761), 
        .A(n6560), .ZN(n6553) );
  AOI221_X1 U4924 ( .B1(net253913), .B2(n37770), .C1(net254105), .C2(n37767), 
        .A(n6559), .ZN(n6554) );
  AOI221_X1 U4925 ( .B1(net253721), .B2(n37776), .C1(net253689), .C2(n37773), 
        .A(n6558), .ZN(n6555) );
  NAND4_X1 U4926 ( .A1(n6511), .A2(n6512), .A3(n6513), .A4(n6514), .ZN(n6510)
         );
  AOI221_X1 U4927 ( .B1(net253594), .B2(n37764), .C1(net253562), .C2(n37761), 
        .A(n6518), .ZN(n6511) );
  AOI221_X1 U4928 ( .B1(net253914), .B2(n37770), .C1(net254106), .C2(n37767), 
        .A(n6517), .ZN(n6512) );
  AOI221_X1 U4929 ( .B1(net253722), .B2(n37776), .C1(net253690), .C2(n37773), 
        .A(n6516), .ZN(n6513) );
  NAND4_X1 U4930 ( .A1(n6341), .A2(n6342), .A3(n6343), .A4(n6344), .ZN(n6340)
         );
  AOI221_X1 U4931 ( .B1(net253595), .B2(n37765), .C1(net253563), .C2(n37762), 
        .A(n6348), .ZN(n6341) );
  AOI221_X1 U4932 ( .B1(net253915), .B2(n37771), .C1(net254107), .C2(n37768), 
        .A(n6347), .ZN(n6342) );
  AOI221_X1 U4933 ( .B1(net253723), .B2(n37777), .C1(net253691), .C2(n37774), 
        .A(n6346), .ZN(n6343) );
  NAND4_X1 U4934 ( .A1(n6299), .A2(n6300), .A3(n6301), .A4(n6302), .ZN(n6298)
         );
  AOI221_X1 U4935 ( .B1(net253596), .B2(n37765), .C1(net253564), .C2(n37762), 
        .A(n6306), .ZN(n6299) );
  AOI221_X1 U4936 ( .B1(net253916), .B2(n37771), .C1(net254108), .C2(n37768), 
        .A(n6305), .ZN(n6300) );
  AOI221_X1 U4937 ( .B1(net253724), .B2(n37777), .C1(net253692), .C2(n37774), 
        .A(n6304), .ZN(n6301) );
  NAND4_X1 U4938 ( .A1(n6257), .A2(n6258), .A3(n6259), .A4(n6260), .ZN(n6256)
         );
  AOI221_X1 U4939 ( .B1(net253597), .B2(n37765), .C1(net253565), .C2(n37762), 
        .A(n6264), .ZN(n6257) );
  AOI221_X1 U4940 ( .B1(net253917), .B2(n37771), .C1(net254109), .C2(n37768), 
        .A(n6263), .ZN(n6258) );
  AOI221_X1 U4941 ( .B1(net253725), .B2(n37777), .C1(net253693), .C2(n37774), 
        .A(n6262), .ZN(n6259) );
  NAND4_X1 U4942 ( .A1(n6215), .A2(n6216), .A3(n6217), .A4(n6218), .ZN(n6214)
         );
  AOI221_X1 U4943 ( .B1(net253598), .B2(n37765), .C1(net253566), .C2(n37762), 
        .A(n6222), .ZN(n6215) );
  AOI221_X1 U4944 ( .B1(net253918), .B2(n37771), .C1(net254110), .C2(n37768), 
        .A(n6221), .ZN(n6216) );
  AOI221_X1 U4945 ( .B1(net253726), .B2(n37777), .C1(net253694), .C2(n37774), 
        .A(n6220), .ZN(n6217) );
  NAND4_X1 U4946 ( .A1(n6173), .A2(n6174), .A3(n6175), .A4(n6176), .ZN(n6172)
         );
  AOI221_X1 U4947 ( .B1(net253599), .B2(n37765), .C1(net253567), .C2(n37762), 
        .A(n6180), .ZN(n6173) );
  AOI221_X1 U4948 ( .B1(net253919), .B2(n37771), .C1(net254111), .C2(n37768), 
        .A(n6179), .ZN(n6174) );
  AOI221_X1 U4949 ( .B1(net253727), .B2(n37777), .C1(net253695), .C2(n37774), 
        .A(n6178), .ZN(n6175) );
  NAND4_X1 U4950 ( .A1(n6131), .A2(n6132), .A3(n6133), .A4(n6134), .ZN(n6130)
         );
  AOI221_X1 U4951 ( .B1(net253600), .B2(n37765), .C1(net253568), .C2(n37762), 
        .A(n6138), .ZN(n6131) );
  AOI221_X1 U4952 ( .B1(net253920), .B2(n37771), .C1(net254112), .C2(n37768), 
        .A(n6137), .ZN(n6132) );
  AOI221_X1 U4953 ( .B1(net253728), .B2(n37777), .C1(net253696), .C2(n37774), 
        .A(n6136), .ZN(n6133) );
  NAND4_X1 U4954 ( .A1(n6089), .A2(n6090), .A3(n6091), .A4(n6092), .ZN(n6088)
         );
  AOI221_X1 U4955 ( .B1(net253601), .B2(n37765), .C1(net253569), .C2(n37762), 
        .A(n6096), .ZN(n6089) );
  AOI221_X1 U4956 ( .B1(net253921), .B2(n37771), .C1(net254113), .C2(n37768), 
        .A(n6095), .ZN(n6090) );
  AOI221_X1 U4957 ( .B1(net253729), .B2(n37777), .C1(net253697), .C2(n37774), 
        .A(n6094), .ZN(n6091) );
  NAND4_X1 U4958 ( .A1(n6047), .A2(n6048), .A3(n6049), .A4(n6050), .ZN(n6046)
         );
  AOI221_X1 U4959 ( .B1(net253602), .B2(n37765), .C1(net253570), .C2(n37762), 
        .A(n6054), .ZN(n6047) );
  AOI221_X1 U4960 ( .B1(net253922), .B2(n37771), .C1(net254114), .C2(n37768), 
        .A(n6053), .ZN(n6048) );
  AOI221_X1 U4961 ( .B1(net253730), .B2(n37777), .C1(net253698), .C2(n37774), 
        .A(n6052), .ZN(n6049) );
  NAND4_X1 U4962 ( .A1(n6005), .A2(n6006), .A3(n6007), .A4(n6008), .ZN(n6004)
         );
  AOI221_X1 U4963 ( .B1(net253603), .B2(n37765), .C1(net253571), .C2(n37762), 
        .A(n6012), .ZN(n6005) );
  AOI221_X1 U4964 ( .B1(net253923), .B2(n37771), .C1(net254115), .C2(n37768), 
        .A(n6011), .ZN(n6006) );
  AOI221_X1 U4965 ( .B1(net253731), .B2(n37777), .C1(net253699), .C2(n37774), 
        .A(n6010), .ZN(n6007) );
  NAND4_X1 U4966 ( .A1(n5963), .A2(n5964), .A3(n5965), .A4(n5966), .ZN(n5962)
         );
  AOI221_X1 U4967 ( .B1(net253604), .B2(n37765), .C1(net253572), .C2(n37762), 
        .A(n5970), .ZN(n5963) );
  AOI221_X1 U4968 ( .B1(net253924), .B2(n37771), .C1(net254116), .C2(n37768), 
        .A(n5969), .ZN(n5964) );
  AOI221_X1 U4969 ( .B1(net253732), .B2(n37777), .C1(net253700), .C2(n37774), 
        .A(n5968), .ZN(n5965) );
  NAND4_X1 U4970 ( .A1(n5921), .A2(n5922), .A3(n5923), .A4(n5924), .ZN(n5920)
         );
  AOI221_X1 U4971 ( .B1(net253605), .B2(n37765), .C1(net253573), .C2(n37762), 
        .A(n5928), .ZN(n5921) );
  AOI221_X1 U4972 ( .B1(net253925), .B2(n37771), .C1(net254117), .C2(n37768), 
        .A(n5927), .ZN(n5922) );
  AOI221_X1 U4973 ( .B1(net253733), .B2(n37777), .C1(net253701), .C2(n37774), 
        .A(n5926), .ZN(n5923) );
  NAND4_X1 U4974 ( .A1(n5879), .A2(n5880), .A3(n5881), .A4(n5882), .ZN(n5878)
         );
  AOI221_X1 U4975 ( .B1(net253606), .B2(n37765), .C1(net253574), .C2(n37762), 
        .A(n5886), .ZN(n5879) );
  AOI221_X1 U4976 ( .B1(net253926), .B2(n37771), .C1(net254118), .C2(n37768), 
        .A(n5885), .ZN(n5880) );
  AOI221_X1 U4977 ( .B1(net253734), .B2(n37777), .C1(net253702), .C2(n37774), 
        .A(n5884), .ZN(n5881) );
  NAND4_X1 U4978 ( .A1(n5837), .A2(n5838), .A3(n5839), .A4(n5840), .ZN(n5836)
         );
  AOI221_X1 U4979 ( .B1(net253607), .B2(n37766), .C1(net253575), .C2(n37763), 
        .A(n5844), .ZN(n5837) );
  AOI221_X1 U4980 ( .B1(net253927), .B2(n37772), .C1(net254119), .C2(n37769), 
        .A(n5843), .ZN(n5838) );
  AOI221_X1 U4981 ( .B1(net253735), .B2(n37778), .C1(net253703), .C2(n37775), 
        .A(n5842), .ZN(n5839) );
  NAND4_X1 U4982 ( .A1(n5795), .A2(n5796), .A3(n5797), .A4(n5798), .ZN(n5794)
         );
  AOI221_X1 U4983 ( .B1(net253608), .B2(n37766), .C1(net253576), .C2(n37763), 
        .A(n5802), .ZN(n5795) );
  AOI221_X1 U4984 ( .B1(net253928), .B2(n37772), .C1(net254120), .C2(n37769), 
        .A(n5801), .ZN(n5796) );
  AOI221_X1 U4985 ( .B1(net253736), .B2(n37778), .C1(net253704), .C2(n37775), 
        .A(n5800), .ZN(n5797) );
  NAND4_X1 U4986 ( .A1(n5753), .A2(n5754), .A3(n5755), .A4(n5756), .ZN(n5752)
         );
  AOI221_X1 U4987 ( .B1(net253609), .B2(n37766), .C1(net253577), .C2(n37763), 
        .A(n5760), .ZN(n5753) );
  AOI221_X1 U4988 ( .B1(net253929), .B2(n37772), .C1(net254121), .C2(n37769), 
        .A(n5759), .ZN(n5754) );
  AOI221_X1 U4989 ( .B1(net253737), .B2(n37778), .C1(net253705), .C2(n37775), 
        .A(n5758), .ZN(n5755) );
  NAND4_X1 U4990 ( .A1(n5711), .A2(n5712), .A3(n5713), .A4(n5714), .ZN(n5710)
         );
  AOI221_X1 U4991 ( .B1(net253610), .B2(n37766), .C1(net253578), .C2(n37763), 
        .A(n5718), .ZN(n5711) );
  AOI221_X1 U4992 ( .B1(net253930), .B2(n37772), .C1(net254122), .C2(n37769), 
        .A(n5717), .ZN(n5712) );
  AOI221_X1 U4993 ( .B1(net253738), .B2(n37778), .C1(net253706), .C2(n37775), 
        .A(n5716), .ZN(n5713) );
  NAND4_X1 U4994 ( .A1(n5669), .A2(n5670), .A3(n5671), .A4(n5672), .ZN(n5668)
         );
  AOI221_X1 U4995 ( .B1(net253611), .B2(n37766), .C1(net253579), .C2(n37763), 
        .A(n5676), .ZN(n5669) );
  AOI221_X1 U4996 ( .B1(net253931), .B2(n37772), .C1(net254123), .C2(n37769), 
        .A(n5675), .ZN(n5670) );
  AOI221_X1 U4997 ( .B1(net253739), .B2(n37778), .C1(net253707), .C2(n37775), 
        .A(n5674), .ZN(n5671) );
  NAND4_X1 U4998 ( .A1(n5627), .A2(n5628), .A3(n5629), .A4(n5630), .ZN(n5626)
         );
  AOI221_X1 U4999 ( .B1(net253612), .B2(n37766), .C1(net253580), .C2(n37763), 
        .A(n5634), .ZN(n5627) );
  AOI221_X1 U5000 ( .B1(net253932), .B2(n37772), .C1(net254124), .C2(n37769), 
        .A(n5633), .ZN(n5628) );
  AOI221_X1 U5001 ( .B1(net253740), .B2(n37778), .C1(net253708), .C2(n37775), 
        .A(n5632), .ZN(n5629) );
  NAND4_X1 U5002 ( .A1(n5585), .A2(n5586), .A3(n5587), .A4(n5588), .ZN(n5584)
         );
  AOI221_X1 U5003 ( .B1(net253613), .B2(n37766), .C1(net253581), .C2(n37763), 
        .A(n5592), .ZN(n5585) );
  AOI221_X1 U5004 ( .B1(net253933), .B2(n37772), .C1(net254125), .C2(n37769), 
        .A(n5591), .ZN(n5586) );
  AOI221_X1 U5005 ( .B1(net253741), .B2(n37778), .C1(net253709), .C2(n37775), 
        .A(n5590), .ZN(n5587) );
  NAND4_X1 U5006 ( .A1(n5518), .A2(n5519), .A3(n5520), .A4(n5521), .ZN(n5517)
         );
  AOI221_X1 U5007 ( .B1(net253614), .B2(n37766), .C1(net253582), .C2(n37763), 
        .A(n5533), .ZN(n5518) );
  AOI221_X1 U5008 ( .B1(net253934), .B2(n37772), .C1(net254126), .C2(n37769), 
        .A(n5530), .ZN(n5519) );
  AOI221_X1 U5009 ( .B1(net253742), .B2(n37778), .C1(net253710), .C2(n37775), 
        .A(n5527), .ZN(n5520) );
  NAND4_X1 U5010 ( .A1(n9592), .A2(n9593), .A3(n9594), .A4(n9595), .ZN(n9564)
         );
  AOI221_X1 U5011 ( .B1(n38557), .B2(n6474), .C1(n38545), .C2(n9613), .A(n9606), .ZN(n9592) );
  AOI221_X1 U5012 ( .B1(n38497), .B2(n6436), .C1(n9609), .C2(n37758), .A(n9600), .ZN(n9593) );
  AOI221_X1 U5013 ( .B1(n38677), .B2(n6402), .C1(n38665), .C2(n9605), .A(n9598), .ZN(n9594) );
  NAND4_X1 U5014 ( .A1(n9531), .A2(n9532), .A3(n9533), .A4(n9534), .ZN(n9521)
         );
  AOI221_X1 U5015 ( .B1(n38557), .B2(n6475), .C1(n38545), .C2(n9548), .A(n9538), .ZN(n9531) );
  AOI221_X1 U5016 ( .B1(n38497), .B2(n6437), .C1(n9546), .C2(n37758), .A(n9537), .ZN(n9532) );
  AOI221_X1 U5017 ( .B1(n38677), .B2(n6403), .C1(n38665), .C2(n9544), .A(n9536), .ZN(n9533) );
  NAND4_X1 U5018 ( .A1(n9489), .A2(n9490), .A3(n9491), .A4(n9492), .ZN(n9479)
         );
  AOI221_X1 U5019 ( .B1(n38557), .B2(n6476), .C1(n38545), .C2(n9506), .A(n9496), .ZN(n9489) );
  AOI221_X1 U5020 ( .B1(n38497), .B2(n6438), .C1(n9504), .C2(n37758), .A(n9495), .ZN(n9490) );
  AOI221_X1 U5021 ( .B1(n38677), .B2(n6404), .C1(n38665), .C2(n9502), .A(n9494), .ZN(n9491) );
  NAND4_X1 U5022 ( .A1(n9447), .A2(n9448), .A3(n9449), .A4(n9450), .ZN(n9437)
         );
  AOI221_X1 U5023 ( .B1(n38557), .B2(n6477), .C1(n38545), .C2(n9464), .A(n9454), .ZN(n9447) );
  AOI221_X1 U5024 ( .B1(n38497), .B2(n6439), .C1(n9462), .C2(n37758), .A(n9453), .ZN(n9448) );
  AOI221_X1 U5025 ( .B1(n38677), .B2(n6405), .C1(n38665), .C2(n9460), .A(n9452), .ZN(n9449) );
  NAND4_X1 U5026 ( .A1(n9405), .A2(n9406), .A3(n9407), .A4(n9408), .ZN(n9395)
         );
  AOI221_X1 U5027 ( .B1(n38557), .B2(n6478), .C1(n38545), .C2(n9422), .A(n9412), .ZN(n9405) );
  AOI221_X1 U5028 ( .B1(n38497), .B2(n6440), .C1(n9420), .C2(n37758), .A(n9411), .ZN(n9406) );
  AOI221_X1 U5029 ( .B1(n38677), .B2(n6407), .C1(n38665), .C2(n9418), .A(n9410), .ZN(n9407) );
  NAND4_X1 U5030 ( .A1(n9363), .A2(n9364), .A3(n9365), .A4(n9366), .ZN(n9353)
         );
  AOI221_X1 U5031 ( .B1(n38557), .B2(n6479), .C1(n38545), .C2(n9380), .A(n9370), .ZN(n9363) );
  AOI221_X1 U5032 ( .B1(n38497), .B2(n6442), .C1(n9378), .C2(n37758), .A(n9369), .ZN(n9364) );
  AOI221_X1 U5033 ( .B1(n38677), .B2(n6409), .C1(n38665), .C2(n9376), .A(n9368), .ZN(n9365) );
  NAND4_X1 U5034 ( .A1(n9321), .A2(n9322), .A3(n9323), .A4(n9324), .ZN(n9311)
         );
  AOI221_X1 U5035 ( .B1(n38557), .B2(n6480), .C1(n38545), .C2(n9338), .A(n9328), .ZN(n9321) );
  AOI221_X1 U5036 ( .B1(n38497), .B2(n6445), .C1(n9336), .C2(n37758), .A(n9327), .ZN(n9322) );
  AOI221_X1 U5037 ( .B1(n38677), .B2(n6410), .C1(n38665), .C2(n9334), .A(n9326), .ZN(n9323) );
  NAND4_X1 U5038 ( .A1(n9279), .A2(n9280), .A3(n9281), .A4(n9282), .ZN(n9269)
         );
  AOI221_X1 U5039 ( .B1(n38557), .B2(n6481), .C1(n38544), .C2(n9296), .A(n9286), .ZN(n9279) );
  AOI221_X1 U5040 ( .B1(n38497), .B2(n6448), .C1(n9294), .C2(n37758), .A(n9285), .ZN(n9280) );
  AOI221_X1 U5041 ( .B1(n38677), .B2(n6411), .C1(n38664), .C2(n9292), .A(n9284), .ZN(n9281) );
  NAND4_X1 U5042 ( .A1(n6645), .A2(n6646), .A3(n6647), .A4(n6648), .ZN(n6635)
         );
  AOI221_X1 U5043 ( .B1(n38557), .B2(n6483), .C1(n38544), .C2(n6662), .A(n6652), .ZN(n6645) );
  AOI221_X1 U5044 ( .B1(n38497), .B2(n6450), .C1(n6660), .C2(n37758), .A(n6651), .ZN(n6646) );
  AOI221_X1 U5045 ( .B1(n38677), .B2(n6412), .C1(n38664), .C2(n6658), .A(n6650), .ZN(n6647) );
  NAND4_X1 U5046 ( .A1(n6603), .A2(n6604), .A3(n6605), .A4(n6606), .ZN(n6593)
         );
  AOI221_X1 U5047 ( .B1(n38556), .B2(n6485), .C1(n38544), .C2(n6620), .A(n6610), .ZN(n6603) );
  AOI221_X1 U5048 ( .B1(n38496), .B2(n6451), .C1(n6618), .C2(n37758), .A(n6609), .ZN(n6604) );
  AOI221_X1 U5049 ( .B1(n38676), .B2(n6413), .C1(n38664), .C2(n6616), .A(n6608), .ZN(n6605) );
  NAND4_X1 U5050 ( .A1(n6561), .A2(n6562), .A3(n6563), .A4(n6564), .ZN(n6551)
         );
  AOI221_X1 U5051 ( .B1(n38556), .B2(n6486), .C1(n38544), .C2(n6578), .A(n6568), .ZN(n6561) );
  AOI221_X1 U5052 ( .B1(n38496), .B2(n6452), .C1(n6576), .C2(n37758), .A(n6567), .ZN(n6562) );
  AOI221_X1 U5053 ( .B1(n38676), .B2(n6414), .C1(n38664), .C2(n6574), .A(n6566), .ZN(n6563) );
  NAND4_X1 U5054 ( .A1(n6519), .A2(n6520), .A3(n6521), .A4(n6522), .ZN(n6509)
         );
  AOI221_X1 U5055 ( .B1(n38556), .B2(n6487), .C1(n38544), .C2(n6536), .A(n6526), .ZN(n6519) );
  AOI221_X1 U5056 ( .B1(n38496), .B2(n6453), .C1(n6534), .C2(n37758), .A(n6525), .ZN(n6520) );
  AOI221_X1 U5057 ( .B1(n38676), .B2(n6415), .C1(n38664), .C2(n6532), .A(n6524), .ZN(n6521) );
  NAND4_X1 U5058 ( .A1(n6349), .A2(n6350), .A3(n6351), .A4(n6352), .ZN(n6339)
         );
  AOI221_X1 U5059 ( .B1(n38556), .B2(n6488), .C1(n38544), .C2(n6366), .A(n6356), .ZN(n6349) );
  AOI221_X1 U5060 ( .B1(n38496), .B2(n6454), .C1(n6364), .C2(n37759), .A(n6355), .ZN(n6350) );
  AOI221_X1 U5061 ( .B1(n38676), .B2(n6416), .C1(n38664), .C2(n6362), .A(n6354), .ZN(n6351) );
  NAND4_X1 U5062 ( .A1(n6307), .A2(n6308), .A3(n6309), .A4(n6310), .ZN(n6297)
         );
  AOI221_X1 U5063 ( .B1(n38556), .B2(n6489), .C1(n38544), .C2(n6324), .A(n6314), .ZN(n6307) );
  AOI221_X1 U5064 ( .B1(n38496), .B2(n6455), .C1(n6322), .C2(n37759), .A(n6313), .ZN(n6308) );
  AOI221_X1 U5065 ( .B1(n38676), .B2(n6417), .C1(n38664), .C2(n6320), .A(n6312), .ZN(n6309) );
  NAND4_X1 U5066 ( .A1(n6265), .A2(n6266), .A3(n6267), .A4(n6268), .ZN(n6255)
         );
  AOI221_X1 U5067 ( .B1(n38556), .B2(n6490), .C1(n38544), .C2(n6282), .A(n6272), .ZN(n6265) );
  AOI221_X1 U5068 ( .B1(n38496), .B2(n6456), .C1(n6280), .C2(n37759), .A(n6271), .ZN(n6266) );
  AOI221_X1 U5069 ( .B1(n38676), .B2(n6418), .C1(n38664), .C2(n6278), .A(n6270), .ZN(n6267) );
  NAND4_X1 U5070 ( .A1(n6223), .A2(n6224), .A3(n6225), .A4(n6226), .ZN(n6213)
         );
  AOI221_X1 U5071 ( .B1(n38556), .B2(n6491), .C1(n38544), .C2(n6240), .A(n6230), .ZN(n6223) );
  AOI221_X1 U5072 ( .B1(n38496), .B2(n6457), .C1(n6238), .C2(n37759), .A(n6229), .ZN(n6224) );
  AOI221_X1 U5073 ( .B1(n38676), .B2(n6419), .C1(n38664), .C2(n6236), .A(n6228), .ZN(n6225) );
  NAND4_X1 U5074 ( .A1(n6181), .A2(n6182), .A3(n6183), .A4(n6184), .ZN(n6171)
         );
  AOI221_X1 U5075 ( .B1(n38556), .B2(n6492), .C1(n38544), .C2(n6198), .A(n6188), .ZN(n6181) );
  AOI221_X1 U5076 ( .B1(n38496), .B2(n6458), .C1(n6196), .C2(n37759), .A(n6187), .ZN(n6182) );
  AOI221_X1 U5077 ( .B1(n38676), .B2(n6420), .C1(n38664), .C2(n6194), .A(n6186), .ZN(n6183) );
  NAND4_X1 U5078 ( .A1(n6139), .A2(n6140), .A3(n6141), .A4(n6142), .ZN(n6129)
         );
  AOI221_X1 U5079 ( .B1(n38556), .B2(n6493), .C1(n38544), .C2(n6156), .A(n6146), .ZN(n6139) );
  AOI221_X1 U5080 ( .B1(n38496), .B2(n6459), .C1(n6154), .C2(n37759), .A(n6145), .ZN(n6140) );
  AOI221_X1 U5081 ( .B1(n38676), .B2(n6421), .C1(n38664), .C2(n6152), .A(n6144), .ZN(n6141) );
  NAND4_X1 U5082 ( .A1(n6097), .A2(n6098), .A3(n6099), .A4(n6100), .ZN(n6087)
         );
  AOI221_X1 U5083 ( .B1(n38556), .B2(n6494), .C1(n38544), .C2(n6114), .A(n6104), .ZN(n6097) );
  AOI221_X1 U5084 ( .B1(n38496), .B2(n6460), .C1(n6112), .C2(n37759), .A(n6103), .ZN(n6098) );
  AOI221_X1 U5085 ( .B1(n38676), .B2(n6422), .C1(n38664), .C2(n6110), .A(n6102), .ZN(n6099) );
  NAND4_X1 U5086 ( .A1(n6055), .A2(n6056), .A3(n6057), .A4(n6058), .ZN(n6045)
         );
  AOI221_X1 U5087 ( .B1(n38556), .B2(n6495), .C1(n38544), .C2(n6072), .A(n6062), .ZN(n6055) );
  AOI221_X1 U5088 ( .B1(n38496), .B2(n6461), .C1(n6070), .C2(n37759), .A(n6061), .ZN(n6056) );
  AOI221_X1 U5089 ( .B1(n38676), .B2(n6423), .C1(n38664), .C2(n6068), .A(n6060), .ZN(n6057) );
  NAND4_X1 U5090 ( .A1(n6013), .A2(n6014), .A3(n6015), .A4(n6016), .ZN(n6003)
         );
  AOI221_X1 U5091 ( .B1(n38556), .B2(n6496), .C1(n38543), .C2(n6030), .A(n6020), .ZN(n6013) );
  AOI221_X1 U5092 ( .B1(n38496), .B2(n6462), .C1(n6028), .C2(n37759), .A(n6019), .ZN(n6014) );
  AOI221_X1 U5093 ( .B1(n38676), .B2(n6424), .C1(n38663), .C2(n6026), .A(n6018), .ZN(n6015) );
  NAND4_X1 U5094 ( .A1(n5971), .A2(n5972), .A3(n5973), .A4(n5974), .ZN(n5961)
         );
  AOI221_X1 U5095 ( .B1(n38555), .B2(n6497), .C1(n38543), .C2(n5988), .A(n5978), .ZN(n5971) );
  AOI221_X1 U5096 ( .B1(n38495), .B2(n6463), .C1(n5986), .C2(n37759), .A(n5977), .ZN(n5972) );
  AOI221_X1 U5097 ( .B1(n38675), .B2(n6425), .C1(n38663), .C2(n5984), .A(n5976), .ZN(n5973) );
  NAND4_X1 U5098 ( .A1(n5929), .A2(n5930), .A3(n5931), .A4(n5932), .ZN(n5919)
         );
  AOI221_X1 U5099 ( .B1(n38555), .B2(n6498), .C1(n38543), .C2(n5946), .A(n5936), .ZN(n5929) );
  AOI221_X1 U5100 ( .B1(n38495), .B2(n6464), .C1(n5944), .C2(n37759), .A(n5935), .ZN(n5930) );
  AOI221_X1 U5101 ( .B1(n38675), .B2(n6426), .C1(n38663), .C2(n5942), .A(n5934), .ZN(n5931) );
  NAND4_X1 U5102 ( .A1(n5887), .A2(n5888), .A3(n5889), .A4(n5890), .ZN(n5877)
         );
  AOI221_X1 U5103 ( .B1(n38555), .B2(n6499), .C1(n38543), .C2(n5904), .A(n5894), .ZN(n5887) );
  AOI221_X1 U5104 ( .B1(n38495), .B2(n6465), .C1(n5902), .C2(n37759), .A(n5893), .ZN(n5888) );
  AOI221_X1 U5105 ( .B1(n38675), .B2(n6427), .C1(n38663), .C2(n5900), .A(n5892), .ZN(n5889) );
  NAND4_X1 U5106 ( .A1(n5845), .A2(n5846), .A3(n5847), .A4(n5848), .ZN(n5835)
         );
  AOI221_X1 U5107 ( .B1(n38555), .B2(n6500), .C1(n38543), .C2(n5862), .A(n5852), .ZN(n5845) );
  AOI221_X1 U5108 ( .B1(n38495), .B2(n6466), .C1(n5860), .C2(n37760), .A(n5851), .ZN(n5846) );
  AOI221_X1 U5109 ( .B1(n38675), .B2(n6428), .C1(n38663), .C2(n5858), .A(n5850), .ZN(n5847) );
  NAND4_X1 U5110 ( .A1(n5803), .A2(n5804), .A3(n5805), .A4(n5806), .ZN(n5793)
         );
  AOI221_X1 U5111 ( .B1(n38555), .B2(n6501), .C1(n38543), .C2(n5820), .A(n5810), .ZN(n5803) );
  AOI221_X1 U5112 ( .B1(n38495), .B2(n6467), .C1(n5818), .C2(n37760), .A(n5809), .ZN(n5804) );
  AOI221_X1 U5113 ( .B1(n38675), .B2(n6429), .C1(n38663), .C2(n5816), .A(n5808), .ZN(n5805) );
  NAND4_X1 U5114 ( .A1(n5761), .A2(n5762), .A3(n5763), .A4(n5764), .ZN(n5751)
         );
  AOI221_X1 U5115 ( .B1(n38555), .B2(n6502), .C1(n38543), .C2(n5778), .A(n5768), .ZN(n5761) );
  AOI221_X1 U5116 ( .B1(n38495), .B2(n6468), .C1(n5776), .C2(n37760), .A(n5767), .ZN(n5762) );
  AOI221_X1 U5117 ( .B1(n38675), .B2(n6430), .C1(n38663), .C2(n5774), .A(n5766), .ZN(n5763) );
  NAND4_X1 U5118 ( .A1(n5719), .A2(n5720), .A3(n5721), .A4(n5722), .ZN(n5709)
         );
  AOI221_X1 U5119 ( .B1(n38555), .B2(n6503), .C1(n38543), .C2(n5736), .A(n5726), .ZN(n5719) );
  AOI221_X1 U5120 ( .B1(n38495), .B2(n6469), .C1(n5734), .C2(n37760), .A(n5725), .ZN(n5720) );
  AOI221_X1 U5121 ( .B1(n38675), .B2(n6431), .C1(n38663), .C2(n5732), .A(n5724), .ZN(n5721) );
  NAND4_X1 U5122 ( .A1(n5677), .A2(n5678), .A3(n5679), .A4(n5680), .ZN(n5667)
         );
  AOI221_X1 U5123 ( .B1(n38555), .B2(n6504), .C1(n38543), .C2(n5694), .A(n5684), .ZN(n5677) );
  AOI221_X1 U5124 ( .B1(n38495), .B2(n6470), .C1(n5692), .C2(n37760), .A(n5683), .ZN(n5678) );
  AOI221_X1 U5125 ( .B1(n38675), .B2(n6432), .C1(n38663), .C2(n5690), .A(n5682), .ZN(n5679) );
  NAND4_X1 U5126 ( .A1(n5635), .A2(n5636), .A3(n5637), .A4(n5638), .ZN(n5625)
         );
  AOI221_X1 U5127 ( .B1(n38555), .B2(n6505), .C1(n38543), .C2(n5652), .A(n5642), .ZN(n5635) );
  AOI221_X1 U5128 ( .B1(n38495), .B2(n6471), .C1(n5650), .C2(n37760), .A(n5641), .ZN(n5636) );
  AOI221_X1 U5129 ( .B1(n38675), .B2(n6433), .C1(n38663), .C2(n5648), .A(n5640), .ZN(n5637) );
  NAND4_X1 U5130 ( .A1(n5593), .A2(n5594), .A3(n5595), .A4(n5596), .ZN(n5583)
         );
  AOI221_X1 U5131 ( .B1(n38555), .B2(n6506), .C1(n38543), .C2(n5610), .A(n5600), .ZN(n5593) );
  AOI221_X1 U5132 ( .B1(n38495), .B2(n6472), .C1(n5608), .C2(n37760), .A(n5599), .ZN(n5594) );
  AOI221_X1 U5133 ( .B1(n38675), .B2(n6434), .C1(n38663), .C2(n5606), .A(n5598), .ZN(n5595) );
  NAND4_X1 U5134 ( .A1(n5534), .A2(n5535), .A3(n5536), .A4(n5537), .ZN(n5516)
         );
  AOI221_X1 U5135 ( .B1(n38555), .B2(n6507), .C1(n38543), .C2(n5560), .A(n5542), .ZN(n5534) );
  AOI221_X1 U5136 ( .B1(n38495), .B2(n6473), .C1(n5558), .C2(n37760), .A(n5541), .ZN(n5535) );
  AOI221_X1 U5137 ( .B1(n38675), .B2(n6435), .C1(n38663), .C2(n5555), .A(n5539), .ZN(n5536) );
  NAND2_X1 U5138 ( .A1(DATAIN[0]), .A2(n38916), .ZN(n2739) );
  NAND2_X1 U5139 ( .A1(DATAIN[1]), .A2(n38916), .ZN(n2737) );
  NAND2_X1 U5140 ( .A1(DATAIN[2]), .A2(n38916), .ZN(n2735) );
  NAND2_X1 U5141 ( .A1(DATAIN[3]), .A2(n38916), .ZN(n2733) );
  NAND2_X1 U5142 ( .A1(DATAIN[4]), .A2(n38916), .ZN(n2731) );
  NAND2_X1 U5143 ( .A1(DATAIN[5]), .A2(n38916), .ZN(n2729) );
  NAND2_X1 U5144 ( .A1(DATAIN[6]), .A2(n38916), .ZN(n2727) );
  NAND2_X1 U5145 ( .A1(DATAIN[7]), .A2(n38916), .ZN(n2725) );
  NAND2_X1 U5146 ( .A1(DATAIN[8]), .A2(n38916), .ZN(n2723) );
  NAND2_X1 U5147 ( .A1(DATAIN[9]), .A2(n38916), .ZN(n2721) );
  NAND2_X1 U5148 ( .A1(DATAIN[10]), .A2(n38916), .ZN(n2719) );
  NAND2_X1 U5149 ( .A1(DATAIN[11]), .A2(n38916), .ZN(n2717) );
  NAND2_X1 U5150 ( .A1(DATAIN[12]), .A2(n38919), .ZN(n2715) );
  NAND2_X1 U5151 ( .A1(DATAIN[13]), .A2(n38918), .ZN(n2713) );
  NAND2_X1 U5152 ( .A1(DATAIN[14]), .A2(n38920), .ZN(n2711) );
  NAND2_X1 U5153 ( .A1(DATAIN[15]), .A2(n38917), .ZN(n2709) );
  NAND2_X1 U5154 ( .A1(DATAIN[16]), .A2(n38916), .ZN(n2707) );
  NAND2_X1 U5155 ( .A1(DATAIN[17]), .A2(n38916), .ZN(n2705) );
  NAND2_X1 U5156 ( .A1(DATAIN[18]), .A2(n38916), .ZN(n2703) );
  NAND2_X1 U5157 ( .A1(DATAIN[19]), .A2(n38916), .ZN(n2701) );
  NAND2_X1 U5158 ( .A1(DATAIN[20]), .A2(n38916), .ZN(n2699) );
  NAND2_X1 U5159 ( .A1(DATAIN[21]), .A2(n38916), .ZN(n2697) );
  NAND2_X1 U5160 ( .A1(DATAIN[22]), .A2(n38920), .ZN(n2695) );
  NAND2_X1 U5161 ( .A1(DATAIN[23]), .A2(n38916), .ZN(n2693) );
  NAND2_X1 U5162 ( .A1(DATAIN[24]), .A2(n38917), .ZN(n2691) );
  NAND2_X1 U5163 ( .A1(DATAIN[25]), .A2(n38919), .ZN(n2689) );
  NAND2_X1 U5164 ( .A1(DATAIN[26]), .A2(n38916), .ZN(n2687) );
  NAND2_X1 U5165 ( .A1(DATAIN[27]), .A2(n38920), .ZN(n2685) );
  NAND2_X1 U5166 ( .A1(DATAIN[28]), .A2(n38919), .ZN(n2683) );
  NAND2_X1 U5167 ( .A1(DATAIN[29]), .A2(n38917), .ZN(n2681) );
  NAND2_X1 U5168 ( .A1(DATAIN[30]), .A2(n38916), .ZN(n2679) );
  NAND2_X1 U5169 ( .A1(DATAIN[31]), .A2(n38920), .ZN(n2677) );
  OR2_X1 U5170 ( .A1(n2812), .A2(Addr[6]), .ZN(n3303) );
  BUF_X1 U5171 ( .A(RESET), .Z(n38914) );
  BUF_X1 U5172 ( .A(RESET), .Z(n38915) );
  NOR2_X1 U5173 ( .A1(n9614), .A2(Addr[3]), .ZN(n9625) );
  AND3_X1 U5174 ( .A1(n9601), .A2(n9604), .A3(Addr[1]), .ZN(n9584) );
  AND3_X1 U5175 ( .A1(Addr[0]), .A2(n9601), .A3(Addr[1]), .ZN(n9599) );
  AND3_X1 U5176 ( .A1(Addr[1]), .A2(Addr[0]), .A3(n9625), .ZN(n9577) );
  AND3_X1 U5177 ( .A1(Addr[2]), .A2(n9604), .A3(n9615), .ZN(n9591) );
  AND3_X1 U5178 ( .A1(Addr[2]), .A2(n9604), .A3(n9619), .ZN(n9571) );
  AND3_X1 U5179 ( .A1(Addr[0]), .A2(n9614), .A3(n9619), .ZN(n9575) );
  AND3_X1 U5180 ( .A1(Addr[2]), .A2(Addr[0]), .A3(n9619), .ZN(n9572) );
  NOR2_X1 U5181 ( .A1(Addr[2]), .A2(Addr[3]), .ZN(n9601) );
  AND3_X1 U5182 ( .A1(n9601), .A2(n9603), .A3(Addr[0]), .ZN(n9587) );
  AND3_X1 U5183 ( .A1(Addr[0]), .A2(n9603), .A3(n9625), .ZN(n9580) );
  AND3_X1 U5184 ( .A1(Addr[1]), .A2(n9604), .A3(n9625), .ZN(n9579) );
  AND3_X1 U5185 ( .A1(Addr[0]), .A2(n9614), .A3(n9615), .ZN(n9573) );
  AND3_X1 U5186 ( .A1(Addr[2]), .A2(Addr[0]), .A3(n9615), .ZN(n9590) );
  INV_X1 U5187 ( .A(Addr[0]), .ZN(n9604) );
  INV_X1 U5188 ( .A(Addr[5]), .ZN(n9630) );
  INV_X1 U5189 ( .A(Addr[4]), .ZN(n9629) );
  INV_X1 U5190 ( .A(Addr[2]), .ZN(n9614) );
  NAND2_X1 U5191 ( .A1(Addr[6]), .A2(n9571), .ZN(n5437) );
  NAND2_X1 U5192 ( .A1(Addr[6]), .A2(n9572), .ZN(n5472) );
  NAND2_X1 U5193 ( .A1(Addr[6]), .A2(n9577), .ZN(n5262) );
  NAND2_X1 U5194 ( .A1(Addr[6]), .A2(n9578), .ZN(n5297) );
  NAND2_X1 U5195 ( .A1(Addr[6]), .A2(n9584), .ZN(n5087) );
  NAND2_X1 U5196 ( .A1(Addr[6]), .A2(n9599), .ZN(n5122) );
  NAND2_X1 U5197 ( .A1(Addr[6]), .A2(n9573), .ZN(n5402) );
  NAND2_X1 U5198 ( .A1(Addr[6]), .A2(n9579), .ZN(n5227) );
  NAND2_X1 U5199 ( .A1(Addr[6]), .A2(n9587), .ZN(n5052) );
  INV_X1 U5200 ( .A(Addr[1]), .ZN(n9603) );
  NAND2_X1 U5201 ( .A1(Addr[6]), .A2(n9575), .ZN(n5332) );
  NAND2_X1 U5202 ( .A1(Addr[6]), .A2(n9581), .ZN(n5157) );
  NAND2_X1 U5203 ( .A1(Addr[6]), .A2(n9591), .ZN(n5507) );
  NAND2_X1 U5204 ( .A1(Addr[6]), .A2(n9574), .ZN(n5367) );
  NAND2_X1 U5205 ( .A1(Addr[6]), .A2(n9580), .ZN(n5192) );
  NAND2_X1 U5206 ( .A1(Addr[6]), .A2(n9590), .ZN(n9560) );
  NAND2_X1 U5207 ( .A1(Addr[6]), .A2(n9589), .ZN(n5017) );
  AND2_X1 U5208 ( .A1(Addr[3]), .A2(n9603), .ZN(n9619) );
  AND2_X1 U5209 ( .A1(Addr[3]), .A2(Addr[1]), .ZN(n9615) );
  CLKBUF_X1 U5210 ( .A(n2739), .Z(n38684) );
  CLKBUF_X1 U5211 ( .A(n2737), .Z(n38691) );
  CLKBUF_X1 U5212 ( .A(n2735), .Z(n38698) );
  CLKBUF_X1 U5213 ( .A(n2733), .Z(n38705) );
  CLKBUF_X1 U5214 ( .A(n2731), .Z(n38712) );
  CLKBUF_X1 U5215 ( .A(n2729), .Z(n38719) );
  CLKBUF_X1 U5216 ( .A(n2727), .Z(n38726) );
  CLKBUF_X1 U5217 ( .A(n2725), .Z(n38733) );
  CLKBUF_X1 U5218 ( .A(n2723), .Z(n38740) );
  CLKBUF_X1 U5219 ( .A(n2721), .Z(n38747) );
  CLKBUF_X1 U5220 ( .A(n2719), .Z(n38754) );
  CLKBUF_X1 U5221 ( .A(n2717), .Z(n38761) );
  CLKBUF_X1 U5222 ( .A(n2715), .Z(n38768) );
  CLKBUF_X1 U5223 ( .A(n2713), .Z(n38775) );
  CLKBUF_X1 U5224 ( .A(n2711), .Z(n38782) );
  CLKBUF_X1 U5225 ( .A(n2709), .Z(n38789) );
  CLKBUF_X1 U5226 ( .A(n2707), .Z(n38796) );
  CLKBUF_X1 U5227 ( .A(n2705), .Z(n38803) );
  CLKBUF_X1 U5228 ( .A(n2703), .Z(n38810) );
  CLKBUF_X1 U5229 ( .A(n2701), .Z(n38817) );
  CLKBUF_X1 U5230 ( .A(n2699), .Z(n38824) );
  CLKBUF_X1 U5231 ( .A(n2697), .Z(n38831) );
  CLKBUF_X1 U5232 ( .A(n2695), .Z(n38838) );
  CLKBUF_X1 U5233 ( .A(n2693), .Z(n38845) );
  CLKBUF_X1 U5234 ( .A(n2691), .Z(n38852) );
  CLKBUF_X1 U5235 ( .A(n2689), .Z(n38859) );
  CLKBUF_X1 U5236 ( .A(n2687), .Z(n38866) );
  CLKBUF_X1 U5237 ( .A(n2685), .Z(n38873) );
  CLKBUF_X1 U5238 ( .A(n2683), .Z(n38880) );
  CLKBUF_X1 U5239 ( .A(n2681), .Z(n38887) );
  CLKBUF_X1 U5240 ( .A(n2679), .Z(n38894) );
  CLKBUF_X1 U5241 ( .A(n2677), .Z(n38901) );
endmodule


module MUX51_GENERIC_N32 ( A, B, C, D, E, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246;

  BUF_X1 U1 ( .A(n240), .Z(n241) );
  BUF_X1 U2 ( .A(n240), .Z(n242) );
  BUF_X1 U3 ( .A(n240), .Z(n243) );
  BUF_X1 U4 ( .A(n6), .Z(n240) );
  NOR4_X1 U5 ( .A1(n237), .A2(n244), .A3(n234), .A4(n231), .ZN(n6) );
  BUF_X1 U6 ( .A(n9), .Z(n232) );
  BUF_X1 U7 ( .A(n8), .Z(n236) );
  BUF_X1 U8 ( .A(n5), .Z(n244) );
  BUF_X1 U9 ( .A(n5), .Z(n245) );
  BUF_X1 U10 ( .A(n8), .Z(n234) );
  BUF_X1 U11 ( .A(n8), .Z(n235) );
  BUF_X1 U12 ( .A(n9), .Z(n231) );
  BUF_X1 U13 ( .A(n7), .Z(n239) );
  BUF_X1 U14 ( .A(n7), .Z(n237) );
  BUF_X1 U15 ( .A(n7), .Z(n238) );
  BUF_X1 U16 ( .A(n9), .Z(n233) );
  BUF_X1 U17 ( .A(n5), .Z(n246) );
  NOR3_X1 U18 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n72), .ZN(n8) );
  NOR3_X1 U19 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n9) );
  AND3_X1 U20 ( .A1(SEL[1]), .A2(n73), .A3(SEL[0]), .ZN(n5) );
  AND3_X1 U21 ( .A1(n72), .A2(n73), .A3(SEL[0]), .ZN(n7) );
  INV_X1 U22 ( .A(SEL[1]), .ZN(n72) );
  NAND2_X1 U23 ( .A1(n20), .A2(n21), .ZN(Y[3]) );
  AOI22_X1 U24 ( .A1(C[3]), .A2(n234), .B1(A[3]), .B2(n231), .ZN(n20) );
  AOI222_X1 U25 ( .A1(D[3]), .A2(n246), .B1(E[3]), .B2(n243), .C1(B[3]), .C2(
        n239), .ZN(n21) );
  NAND2_X1 U26 ( .A1(n18), .A2(n19), .ZN(Y[4]) );
  AOI22_X1 U27 ( .A1(C[4]), .A2(n234), .B1(A[4]), .B2(n231), .ZN(n18) );
  AOI222_X1 U28 ( .A1(D[4]), .A2(n246), .B1(E[4]), .B2(n243), .C1(B[4]), .C2(
        n239), .ZN(n19) );
  NAND2_X1 U29 ( .A1(n16), .A2(n17), .ZN(Y[5]) );
  AOI22_X1 U30 ( .A1(C[5]), .A2(n234), .B1(A[5]), .B2(n231), .ZN(n16) );
  AOI222_X1 U31 ( .A1(D[5]), .A2(n246), .B1(E[5]), .B2(n243), .C1(B[5]), .C2(
        n239), .ZN(n17) );
  NAND2_X1 U32 ( .A1(n14), .A2(n15), .ZN(Y[6]) );
  AOI22_X1 U33 ( .A1(C[6]), .A2(n234), .B1(A[6]), .B2(n231), .ZN(n14) );
  AOI222_X1 U34 ( .A1(D[6]), .A2(n246), .B1(E[6]), .B2(n243), .C1(B[6]), .C2(
        n239), .ZN(n15) );
  NAND2_X1 U35 ( .A1(n12), .A2(n13), .ZN(Y[7]) );
  AOI22_X1 U36 ( .A1(C[7]), .A2(n234), .B1(A[7]), .B2(n231), .ZN(n12) );
  AOI222_X1 U37 ( .A1(D[7]), .A2(n246), .B1(E[7]), .B2(n243), .C1(B[7]), .C2(
        n239), .ZN(n13) );
  NAND2_X1 U38 ( .A1(n10), .A2(n11), .ZN(Y[8]) );
  AOI22_X1 U39 ( .A1(C[8]), .A2(n234), .B1(A[8]), .B2(n231), .ZN(n10) );
  AOI222_X1 U40 ( .A1(D[8]), .A2(n246), .B1(E[8]), .B2(n243), .C1(B[8]), .C2(
        n239), .ZN(n11) );
  NAND2_X1 U41 ( .A1(n3), .A2(n4), .ZN(Y[9]) );
  AOI22_X1 U42 ( .A1(C[9]), .A2(n235), .B1(A[9]), .B2(n232), .ZN(n3) );
  AOI222_X1 U43 ( .A1(D[9]), .A2(n246), .B1(E[9]), .B2(n243), .C1(B[9]), .C2(
        n239), .ZN(n4) );
  NAND2_X1 U44 ( .A1(n22), .A2(n23), .ZN(Y[31]) );
  AOI22_X1 U45 ( .A1(C[31]), .A2(n234), .B1(A[31]), .B2(n231), .ZN(n22) );
  AOI222_X1 U46 ( .A1(D[31]), .A2(n245), .B1(E[31]), .B2(n243), .C1(B[31]), 
        .C2(n239), .ZN(n23) );
  NAND2_X1 U47 ( .A1(n24), .A2(n25), .ZN(Y[30]) );
  AOI22_X1 U48 ( .A1(C[30]), .A2(n234), .B1(A[30]), .B2(n231), .ZN(n24) );
  AOI222_X1 U49 ( .A1(D[30]), .A2(n245), .B1(E[30]), .B2(n242), .C1(B[30]), 
        .C2(n239), .ZN(n25) );
  NAND2_X1 U50 ( .A1(n70), .A2(n71), .ZN(Y[0]) );
  AOI22_X1 U51 ( .A1(C[0]), .A2(n234), .B1(A[0]), .B2(n231), .ZN(n70) );
  AOI222_X1 U52 ( .A1(D[0]), .A2(n244), .B1(E[0]), .B2(n241), .C1(B[0]), .C2(
        n237), .ZN(n71) );
  NAND2_X1 U53 ( .A1(n48), .A2(n49), .ZN(Y[1]) );
  AOI22_X1 U54 ( .A1(C[1]), .A2(n235), .B1(A[1]), .B2(n232), .ZN(n48) );
  AOI222_X1 U55 ( .A1(D[1]), .A2(n244), .B1(E[1]), .B2(n241), .C1(B[1]), .C2(
        n238), .ZN(n49) );
  NAND2_X1 U56 ( .A1(n26), .A2(n27), .ZN(Y[2]) );
  AOI22_X1 U57 ( .A1(C[2]), .A2(n234), .B1(A[2]), .B2(n231), .ZN(n26) );
  AOI222_X1 U58 ( .A1(D[2]), .A2(n245), .B1(E[2]), .B2(n242), .C1(B[2]), .C2(
        n238), .ZN(n27) );
  NAND2_X1 U59 ( .A1(n68), .A2(n69), .ZN(Y[10]) );
  AOI22_X1 U60 ( .A1(C[10]), .A2(n236), .B1(A[10]), .B2(n233), .ZN(n68) );
  AOI222_X1 U61 ( .A1(D[10]), .A2(n244), .B1(E[10]), .B2(n241), .C1(B[10]), 
        .C2(n237), .ZN(n69) );
  NAND2_X1 U62 ( .A1(n66), .A2(n67), .ZN(Y[11]) );
  AOI22_X1 U63 ( .A1(C[11]), .A2(n236), .B1(A[11]), .B2(n233), .ZN(n66) );
  AOI222_X1 U64 ( .A1(D[11]), .A2(n244), .B1(E[11]), .B2(n241), .C1(B[11]), 
        .C2(n237), .ZN(n67) );
  NAND2_X1 U65 ( .A1(n64), .A2(n65), .ZN(Y[12]) );
  AOI22_X1 U66 ( .A1(C[12]), .A2(n236), .B1(A[12]), .B2(n233), .ZN(n64) );
  AOI222_X1 U67 ( .A1(D[12]), .A2(n244), .B1(E[12]), .B2(n241), .C1(B[12]), 
        .C2(n237), .ZN(n65) );
  NAND2_X1 U68 ( .A1(n62), .A2(n63), .ZN(Y[13]) );
  AOI22_X1 U69 ( .A1(C[13]), .A2(n236), .B1(A[13]), .B2(n233), .ZN(n62) );
  AOI222_X1 U70 ( .A1(D[13]), .A2(n244), .B1(E[13]), .B2(n241), .C1(B[13]), 
        .C2(n237), .ZN(n63) );
  NAND2_X1 U71 ( .A1(n60), .A2(n61), .ZN(Y[14]) );
  AOI22_X1 U72 ( .A1(C[14]), .A2(n236), .B1(A[14]), .B2(n233), .ZN(n60) );
  AOI222_X1 U73 ( .A1(D[14]), .A2(n244), .B1(E[14]), .B2(n241), .C1(B[14]), 
        .C2(n237), .ZN(n61) );
  NAND2_X1 U74 ( .A1(n58), .A2(n59), .ZN(Y[15]) );
  AOI22_X1 U75 ( .A1(C[15]), .A2(n236), .B1(A[15]), .B2(n233), .ZN(n58) );
  AOI222_X1 U76 ( .A1(D[15]), .A2(n244), .B1(E[15]), .B2(n241), .C1(B[15]), 
        .C2(n237), .ZN(n59) );
  NAND2_X1 U77 ( .A1(n56), .A2(n57), .ZN(Y[16]) );
  AOI22_X1 U78 ( .A1(C[16]), .A2(n236), .B1(A[16]), .B2(n233), .ZN(n56) );
  AOI222_X1 U79 ( .A1(D[16]), .A2(n244), .B1(E[16]), .B2(n241), .C1(B[16]), 
        .C2(n237), .ZN(n57) );
  NAND2_X1 U80 ( .A1(n54), .A2(n55), .ZN(Y[17]) );
  AOI22_X1 U81 ( .A1(C[17]), .A2(n236), .B1(A[17]), .B2(n233), .ZN(n54) );
  AOI222_X1 U82 ( .A1(D[17]), .A2(n244), .B1(E[17]), .B2(n241), .C1(B[17]), 
        .C2(n237), .ZN(n55) );
  NAND2_X1 U83 ( .A1(n52), .A2(n53), .ZN(Y[18]) );
  AOI22_X1 U84 ( .A1(C[18]), .A2(n236), .B1(A[18]), .B2(n232), .ZN(n52) );
  AOI222_X1 U85 ( .A1(D[18]), .A2(n244), .B1(E[18]), .B2(n241), .C1(B[18]), 
        .C2(n237), .ZN(n53) );
  NAND2_X1 U86 ( .A1(n50), .A2(n51), .ZN(Y[19]) );
  AOI22_X1 U87 ( .A1(C[19]), .A2(n235), .B1(A[19]), .B2(n232), .ZN(n50) );
  AOI222_X1 U88 ( .A1(D[19]), .A2(n244), .B1(E[19]), .B2(n241), .C1(B[19]), 
        .C2(n237), .ZN(n51) );
  NAND2_X1 U89 ( .A1(n46), .A2(n47), .ZN(Y[20]) );
  AOI22_X1 U90 ( .A1(C[20]), .A2(n235), .B1(A[20]), .B2(n232), .ZN(n46) );
  AOI222_X1 U91 ( .A1(D[20]), .A2(n245), .B1(E[20]), .B2(n242), .C1(B[20]), 
        .C2(n238), .ZN(n47) );
  NAND2_X1 U92 ( .A1(n44), .A2(n45), .ZN(Y[21]) );
  AOI22_X1 U93 ( .A1(C[21]), .A2(n235), .B1(A[21]), .B2(n232), .ZN(n44) );
  AOI222_X1 U94 ( .A1(D[21]), .A2(n245), .B1(E[21]), .B2(n242), .C1(B[21]), 
        .C2(n238), .ZN(n45) );
  NAND2_X1 U95 ( .A1(n42), .A2(n43), .ZN(Y[22]) );
  AOI22_X1 U96 ( .A1(C[22]), .A2(n235), .B1(A[22]), .B2(n232), .ZN(n42) );
  AOI222_X1 U97 ( .A1(D[22]), .A2(n245), .B1(E[22]), .B2(n242), .C1(B[22]), 
        .C2(n238), .ZN(n43) );
  NAND2_X1 U98 ( .A1(n40), .A2(n41), .ZN(Y[23]) );
  AOI22_X1 U99 ( .A1(C[23]), .A2(n235), .B1(A[23]), .B2(n232), .ZN(n40) );
  AOI222_X1 U100 ( .A1(D[23]), .A2(n245), .B1(E[23]), .B2(n242), .C1(B[23]), 
        .C2(n238), .ZN(n41) );
  NAND2_X1 U101 ( .A1(n38), .A2(n39), .ZN(Y[24]) );
  AOI22_X1 U102 ( .A1(C[24]), .A2(n235), .B1(A[24]), .B2(n232), .ZN(n38) );
  AOI222_X1 U103 ( .A1(D[24]), .A2(n245), .B1(E[24]), .B2(n242), .C1(B[24]), 
        .C2(n238), .ZN(n39) );
  NAND2_X1 U104 ( .A1(n36), .A2(n37), .ZN(Y[25]) );
  AOI22_X1 U105 ( .A1(C[25]), .A2(n235), .B1(A[25]), .B2(n232), .ZN(n36) );
  AOI222_X1 U106 ( .A1(D[25]), .A2(n245), .B1(E[25]), .B2(n242), .C1(B[25]), 
        .C2(n238), .ZN(n37) );
  NAND2_X1 U107 ( .A1(n34), .A2(n35), .ZN(Y[26]) );
  AOI22_X1 U108 ( .A1(C[26]), .A2(n235), .B1(A[26]), .B2(n232), .ZN(n34) );
  AOI222_X1 U109 ( .A1(D[26]), .A2(n245), .B1(E[26]), .B2(n242), .C1(B[26]), 
        .C2(n238), .ZN(n35) );
  NAND2_X1 U110 ( .A1(n32), .A2(n33), .ZN(Y[27]) );
  AOI22_X1 U111 ( .A1(C[27]), .A2(n235), .B1(A[27]), .B2(n232), .ZN(n32) );
  AOI222_X1 U112 ( .A1(D[27]), .A2(n245), .B1(E[27]), .B2(n242), .C1(B[27]), 
        .C2(n238), .ZN(n33) );
  NAND2_X1 U113 ( .A1(n30), .A2(n31), .ZN(Y[28]) );
  AOI22_X1 U114 ( .A1(C[28]), .A2(n235), .B1(A[28]), .B2(n232), .ZN(n30) );
  AOI222_X1 U115 ( .A1(D[28]), .A2(n245), .B1(E[28]), .B2(n242), .C1(B[28]), 
        .C2(n238), .ZN(n31) );
  NAND2_X1 U116 ( .A1(n28), .A2(n29), .ZN(Y[29]) );
  AOI22_X1 U117 ( .A1(C[29]), .A2(n234), .B1(A[29]), .B2(n231), .ZN(n28) );
  AOI222_X1 U118 ( .A1(D[29]), .A2(n245), .B1(E[29]), .B2(n242), .C1(B[29]), 
        .C2(n238), .ZN(n29) );
  INV_X1 U119 ( .A(SEL[2]), .ZN(n73) );
endmodule


module ALU_N32 ( ALU_OPCODE, A, B, Y_ADDER, Y_SHIFT, Y_LOGIC, Y_MULT, ne, ge, 
        le, ee );
  input [7:0] ALU_OPCODE;
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y_ADDER;
  output [31:0] Y_SHIFT;
  output [31:0] Y_LOGIC;
  output [31:0] Y_MULT;
  output ne, ge, le, ee;
  wire   carry, n1, n2, n3, n4, n5, n6, n7, n8, n9, n11, n12, n13, n14, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n34, n35;
  assign n1 = B[7];
  assign n2 = B[4];
  assign n3 = A[4];
  assign n4 = B[2];
  assign n5 = A[6];
  assign n6 = A[12];
  assign n7 = A[14];
  assign n8 = B[0];
  assign n9 = B[3];
  assign n11 = A[0];
  assign n12 = A[1];
  assign n13 = A[2];
  assign n14 = A[3];
  assign n16 = A[5];
  assign n17 = A[7];
  assign n18 = A[8];
  assign n19 = A[9];
  assign n20 = A[10];
  assign n21 = A[11];
  assign n22 = A[13];
  assign n23 = A[15];
  assign n24 = A[16];
  assign n25 = A[18];
  assign n26 = A[20];
  assign n27 = A[22];
  assign n34 = B[1];

  Logic_Unit_N32 Logic_unit_exe ( .R1({A[31:23], n27, A[21], n26, A[19], n25, 
        A[17], n24, n23, n7, n22, n6, n21, n20, n19, n18, n17, n5, n16, n3, 
        n14, n13, n12, n11}), .R2({B[31:8], n1, B[6:5], n2, n9, n4, n35, n8}), 
        .S1(ALU_OPCODE[2]), .S2(ALU_OPCODE[1]), .S3(ALU_OPCODE[0]), .S0(
        ALU_OPCODE[3]), .Y(Y_LOGIC) );
  P4adder_subtr_N32_M4 P4Adder_exe ( .A({A[31:23], n27, A[21], n26, A[19], n25, 
        A[17], n24, n23, n7, n22, n6, n21, n20, n19, n18, n17, n5, n16, n3, 
        n14, n13, n12, n11}), .B({B[31:8], n1, B[6:5], n2, n9, n4, n35, n8}), 
        .Y(Y_ADDER), .SEL(ALU_OPCODE[4]), .Co(carry) );
  comparator Comparator_exe ( .SUB(Y_ADDER), .Cout(carry), .ne(ne), .ge(ge), 
        .le(le), .ee(ee) );
  SHIFTER_GENERIC_N32 Shifter_exe ( .A({A[31:23], n27, A[21], n26, A[19], n25, 
        A[17], n24, n23, n7, n22, n6, n21, n20, n19, n18, n17, n5, n16, n3, 
        n14, n13, n12, n11}), .B({n2, n9, n4, n35, n8}), .LOGIC_ARITH(
        ALU_OPCODE[7]), .LEFT_RIGHT(ALU_OPCODE[6]), .SHIFT_ROTATE(
        ALU_OPCODE[5]), .OUTPUT(Y_SHIFT) );
  boothmul_N16_M16 mult_exe ( .Am({n23, n7, n22, n6, n21, n20, n19, n18, n17, 
        n5, n16, n3, n14, n13, n12, n11}), .Bm({B[15:8], n1, B[6:5], n2, n9, 
        n4, n35, n8}), .Pm(Y_MULT) );
  BUF_X1 U1 ( .A(n34), .Z(n35) );
endmodule


module zero_detector_N32 ( A, YE );
  input [31:0] A;
  output YE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  NOR4_X1 U1 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n10) );
  NOR4_X1 U2 ( .A1(A[22]), .A2(A[21]), .A3(A[20]), .A4(A[1]), .ZN(n6) );
  NOR4_X1 U3 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[30]), .ZN(n9) );
  NOR4_X1 U4 ( .A1(A[19]), .A2(A[18]), .A3(A[17]), .A4(A[16]), .ZN(n5) );
  NOR4_X1 U5 ( .A1(A[2]), .A2(A[29]), .A3(A[28]), .A4(A[27]), .ZN(n8) );
  NOR4_X1 U6 ( .A1(A[15]), .A2(A[14]), .A3(A[13]), .A4(A[12]), .ZN(n4) );
  NOR4_X1 U7 ( .A1(A[26]), .A2(A[25]), .A3(A[24]), .A4(A[23]), .ZN(n7) );
  NOR2_X1 U8 ( .A1(n1), .A2(n2), .ZN(YE) );
  NAND4_X1 U9 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(n2) );
  NAND4_X1 U10 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(n1) );
  NOR3_X1 U11 ( .A1(A[0]), .A2(A[11]), .A3(A[10]), .ZN(n3) );
endmodule


module MUX41_GENERIC_N6 ( A, B, C, D, SEL, Y );
  input [5:0] A;
  input [5:0] B;
  input [5:0] C;
  input [5:0] D;
  input [1:0] SEL;
  output [5:0] Y;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18;

  NOR3_X1 U1 ( .A1(n6), .A2(n7), .A3(n5), .ZN(n4) );
  NOR2_X1 U2 ( .A1(n18), .A2(SEL[0]), .ZN(n6) );
  NOR2_X1 U3 ( .A1(SEL[0]), .A2(SEL[1]), .ZN(n7) );
  AND2_X1 U4 ( .A1(SEL[0]), .A2(n18), .ZN(n5) );
  INV_X1 U5 ( .A(SEL[1]), .ZN(n18) );
  NAND2_X1 U6 ( .A1(n16), .A2(n17), .ZN(Y[0]) );
  AOI22_X1 U7 ( .A1(C[0]), .A2(n6), .B1(A[0]), .B2(n7), .ZN(n16) );
  AOI22_X1 U8 ( .A1(D[0]), .A2(n4), .B1(B[0]), .B2(n5), .ZN(n17) );
  NAND2_X1 U9 ( .A1(n14), .A2(n15), .ZN(Y[1]) );
  AOI22_X1 U10 ( .A1(C[1]), .A2(n6), .B1(A[1]), .B2(n7), .ZN(n14) );
  AOI22_X1 U11 ( .A1(D[1]), .A2(n4), .B1(B[1]), .B2(n5), .ZN(n15) );
  NAND2_X1 U12 ( .A1(n12), .A2(n13), .ZN(Y[2]) );
  AOI22_X1 U13 ( .A1(C[2]), .A2(n6), .B1(A[2]), .B2(n7), .ZN(n12) );
  AOI22_X1 U14 ( .A1(D[2]), .A2(n4), .B1(B[2]), .B2(n5), .ZN(n13) );
  NAND2_X1 U15 ( .A1(n10), .A2(n11), .ZN(Y[3]) );
  AOI22_X1 U16 ( .A1(C[3]), .A2(n6), .B1(A[3]), .B2(n7), .ZN(n10) );
  AOI22_X1 U17 ( .A1(D[3]), .A2(n4), .B1(B[3]), .B2(n5), .ZN(n11) );
  NAND2_X1 U18 ( .A1(n8), .A2(n9), .ZN(Y[4]) );
  AOI22_X1 U19 ( .A1(C[4]), .A2(n6), .B1(A[4]), .B2(n7), .ZN(n8) );
  AOI22_X1 U20 ( .A1(D[4]), .A2(n4), .B1(B[4]), .B2(n5), .ZN(n9) );
  NAND2_X1 U21 ( .A1(n2), .A2(n3), .ZN(Y[5]) );
  AOI22_X1 U22 ( .A1(C[5]), .A2(n6), .B1(A[5]), .B2(n7), .ZN(n2) );
  AOI22_X1 U23 ( .A1(D[5]), .A2(n4), .B1(B[5]), .B2(n5), .ZN(n3) );
endmodule


module reg_generic_N5 ( D, CLK, RST, EN, Q );
  input [4:0] D;
  output [4:0] Q;
  input CLK, RST, EN;


  FD_s_261 UFD_0 ( .D(D[0]), .CLK(CLK), .RST(RST), .EN(EN), .Q(Q[0]) );
  FD_s_260 UFD_1 ( .D(D[1]), .CLK(CLK), .RST(RST), .EN(EN), .Q(Q[1]) );
  FD_s_259 UFD_2 ( .D(D[2]), .CLK(CLK), .RST(RST), .EN(EN), .Q(Q[2]) );
  FD_s_258 UFD_3 ( .D(D[3]), .CLK(CLK), .RST(RST), .EN(EN), .Q(Q[3]) );
  FD_s_257 UFD_4 ( .D(D[4]), .CLK(CLK), .RST(RST), .EN(EN), .Q(Q[4]) );
endmodule


module reg_generic_N26 ( D, CLK, RST, EN, Q );
  input [25:0] D;
  output [25:0] Q;
  input CLK, RST, EN;
  wire   n6, n7;
  assign n6 = RST;
  assign n7 = EN;

  FD_s_319 UFD_0 ( .D(D[0]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[0]) );
  FD_s_318 UFD_1 ( .D(D[1]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[1]) );
  FD_s_317 UFD_2 ( .D(D[2]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[2]) );
  FD_s_316 UFD_3 ( .D(D[3]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[3]) );
  FD_s_315 UFD_4 ( .D(D[4]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[4]) );
  FD_s_314 UFD_5 ( .D(D[5]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[5]) );
  FD_s_313 UFD_6 ( .D(D[6]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[6]) );
  FD_s_312 UFD_7 ( .D(D[7]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[7]) );
  FD_s_311 UFD_8 ( .D(D[8]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[8]) );
  FD_s_310 UFD_9 ( .D(D[9]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[9]) );
  FD_s_309 UFD_10 ( .D(D[10]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[10]) );
  FD_s_308 UFD_11 ( .D(D[11]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[11]) );
  FD_s_307 UFD_12 ( .D(D[12]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[12]) );
  FD_s_306 UFD_13 ( .D(D[13]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[13]) );
  FD_s_305 UFD_14 ( .D(D[14]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[14]) );
  FD_s_304 UFD_15 ( .D(D[15]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[15]) );
  FD_s_303 UFD_16 ( .D(D[16]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[16]) );
  FD_s_302 UFD_17 ( .D(D[17]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[17]) );
  FD_s_301 UFD_18 ( .D(D[18]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[18]) );
  FD_s_300 UFD_19 ( .D(D[19]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[19]) );
  FD_s_299 UFD_20 ( .D(D[20]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[20]) );
  FD_s_298 UFD_21 ( .D(D[21]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[21]) );
  FD_s_297 UFD_22 ( .D(D[22]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[22]) );
  FD_s_296 UFD_23 ( .D(D[23]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[23]) );
  FD_s_295 UFD_24 ( .D(D[24]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[24]) );
  FD_s_294 UFD_25 ( .D(D[25]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[25]) );
endmodule


module register_file_N32_A5_tot_regs32 ( CLK, RESET, ENABLE, RD1, RD2, WR, 
        ADD_WR, ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RESET, ENABLE, RD1, RD2, WR;
  wire   n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, net310470,
         net310471, net310472, net310473, net310474, net310475, net310476,
         net310477, net310478, net310479, net310480, net310481, net310482,
         net310483, net310484, net310485, net310486, net310487, net310488,
         net310489, net310490, net310491, net310492, net310493, net310494,
         net310495, net310496, net310497, net310498, net310499, net310500,
         net310502, net310503, net310504, net310505, net310506, net310507,
         net310508, net310509, net310510, net310511, net310512, net310513,
         net310514, net310515, net310516, net310517, net310518, net310519,
         net310520, net310521, net310522, net310523, net310524, net310525,
         net310526, net310527, net310528, net310529, net310530, net310531,
         net310532, net310533, net310758, net310759, net310760, net310761,
         net310762, net310763, net310764, net310765, net310766, net310767,
         net310768, net310769, net310770, net310771, net310772, net310773,
         net310774, net310775, net310776, net310777, net310778, net310779,
         net310780, net310781, net310782, net310783, net310784, net310785,
         net310786, net310787, net310788, net310789, net366951, net366952,
         net366953, net366954, net366955, net366956, net366957, net366958,
         net366959, net366960, net366961, net366962, net366963, net366964,
         net366965, net366966, net366967, net366968, net366969, net366970,
         net366971, net366972, net366973, net366974, net366975, net366976,
         net366977, net366978, net366979, net366980, net366981, net366982,
         net367015, net367016, net367017, net367018, net367019, net367020,
         net367021, net367022, net367023, net367024, net367025, net367026,
         net367027, net367028, net367029, net367030, net367031, net367032,
         net367033, net367034, net367035, net367036, net367037, net367038,
         net367039, net367040, net367041, net367042, net367043, net367044,
         net367045, net367046, net367111, net367112, net367113, net367114,
         net367115, net367116, net367117, net367118, net367119, net367120,
         net367121, net367122, net367123, net367124, net367125, net367126,
         net367127, net367128, net367129, net367130, net367131, net367132,
         net367133, net367134, net367135, net367136, net367137, net367138,
         net367139, net367140, net367141, net367142, net423174, net423175,
         net423176, net423177, net423178, net423179, net423180, net423181,
         net423182, net423183, net423184, net423185, net423186, net423187,
         net423188, net423189, net423190, net423191, net423192, net423193,
         net423194, net423195, net423196, net423197, net423198, net423199,
         net423200, net423201, net423202, net423203, net423204, net423205,
         net423334, net423335, net423336, net423337, net423338, net423339,
         net423340, net423341, net423342, net423343, net423344, net423345,
         net423346, net423347, net423348, net423349, net423350, net423351,
         net423352, net423353, net423354, net423355, net423356, net423357,
         net423358, net423359, net423360, net423361, net423362, net423363,
         net423364, net423365, net479344, net479345, net479346, net479347,
         net479348, net479349, net479350, net479351, net479352, net479353,
         net479354, net479355, net479356, net479357, net479358, net479359,
         net479360, net479361, net479362, net479363, net479364, net479365,
         net479366, net479367, net479368, net479369, net479370, net479371,
         net479372, net479373, net479374, net479375, net479376, net479377,
         net479378, net479379, net479380, net479381, net479382, net479383,
         net479384, net479385, net479386, net479387, net479388, net479389,
         net479390, net479391, net479392, net479393, net479394, net479395,
         net479396, net479397, net479398, net479399, net479400, net479401,
         net479402, net479403, net479404, net479405, net479406, net479407,
         net479408, net479410, net479411, net479412, net479413, net479414,
         net479415, net479416, net479417, net479418, net479419, net479420,
         net479421, net479422, net479423, net479424, net479425, net479426,
         net479427, net479428, net479429, net479430, net479431, net479432,
         net479433, net479434, net479435, net479436, net479437, net479438,
         net479439, net479440, net479441, net535436, net535437, net535438,
         net535439, net535440, net535441, net535442, net535443, net535444,
         net535445, net535446, net535447, net535448, net535449, net535450,
         net535451, net535452, net535453, net535454, net535455, net535456,
         net535457, net535458, net535459, net535460, net535461, net535462,
         net535463, net535464, net535465, net535466, net535467, net535468,
         net535469, net535470, net535471, net535472, net535473, net535474,
         net535475, net535476, net535477, net535478, net535479, net535480,
         net535481, net535482, net535483, net535484, net535485, net535486,
         net535487, net535488, net535489, net535490, net535491, net535492,
         net535493, net535494, net535495, net535496, net535497, net535498,
         net535499, net535500, net535501, net535502, net535503, net535504,
         net535505, net535506, net535507, net535508, net535509, net535510,
         net535511, net535512, net535513, net535514, net535515, net535516,
         net535517, net535518, net535519, net535520, net535521, net535522,
         net535523, net535524, net535525, net535526, net535527, net535528,
         net535529, net535530, net535531, net535532, net535533, net535534,
         net535535, net535536, net535537, net535538, net535539, net535540,
         net535541, net535542, net535543, net535544, net535545, net535546,
         net535547, net535548, net535549, net535550, net535551, net535552,
         net535553, net535554, net535555, net535556, net535557, net535558,
         net535559, net535560, net535561, net535562, net535563, net591531,
         net591532, net591533, net591534, net591535, net591536, net591537,
         net591538, net591539, net591540, net591541, net591542, net591543,
         net591544, net591545, net591546, net591547, net591548, net591549,
         net591550, net591551, net591552, net591553, net591554, net591555,
         net591556, net591557, net591558, net591559, net591560, net591561,
         net591562, net591627, net591628, net591629, net591630, net591631,
         net591632, net591633, net591634, net591635, net591636, net591637,
         net591638, net591639, net591640, net591641, net591642, net591643,
         net591644, net591645, net591646, net591647, net591648, net591649,
         net591650, net591651, net591652, net591653, net591654, net591655,
         net591656, net591657, net591658, net591659, net591660, net591661,
         net591662, net591663, net591664, net591665, net591666, net591667,
         net591668, net591669, net591670, net591671, net591672, net591673,
         net591674, net591675, net591676, net591677, net591678, net591679,
         net591680, net591681, net591682, net591683, net591684, net591685,
         net591686, net591687, net591688, net591689, net591690, net591723,
         net591724, net591725, net591726, net591727, net591728, net591729,
         net591730, net591731, net591732, net591733, net591734, net591735,
         net591736, net591737, net591738, net591739, net591740, net591741,
         net591742, net591743, net591744, net591745, net591746, net591747,
         net591748, net591749, net591750, net591751, net591752, net591753,
         net591754, net591787, net591788, net591789, net591790, net591791,
         net591792, net591793, net591794, net591795, net591796, net591797,
         net591798, net591799, net591800, net591801, net591802, net591803,
         net591804, net591805, net591806, net591807, net591808, net591809,
         net591810, net591811, net591812, net591813, net591814, net591815,
         net591816, net591817, net591818, n1073, n1074, n1076, n1078, n1080,
         n1082, n1084, n1086, n1088, n1090, n1092, n1094, n1096, n1098, n1100,
         n1102, n1104, n1106, n1108, n1110, n1112, n1114, n1116, n1118, n1120,
         n1122, n1124, n1126, n1128, n1130, n1132, n1134, n1136, n1138, n1139,
         n1142, n1174, n1176, n1178, n1209, n1212, n1214, n1247, n1248, n1249,
         n1250, n1252, n1282, n1286, n1288, n1322, n1356, n1390, n1419, n1424,
         n1426, n1460, n1494, n1528, n1561, n1563, n1597, n1631, n1664, n1666,
         n1694, n1700, n1702, n1736, n1770, n1803, n1805, n1838, n1840, n1874,
         n1908, n1942, n1975, n1977, n2011, n2045, n2079, n2112, n2113, n2114,
         n2116, n2150, n2183, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4553, n4554, n4555,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
         n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
         n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
         n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686,
         n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
         n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
         n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
         n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
         n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
         n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
         n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
         n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
         n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
         n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798,
         n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
         n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
         n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
         n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830,
         n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
         n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
         n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
         n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
         n18999;

  DFF_X1 \REGISTERS_reg[0][31]  ( .D(n3847), .CK(CLK), .Q(net310789), .QN(
        n17943) );
  DFF_X1 \REGISTERS_reg[0][30]  ( .D(n3846), .CK(CLK), .Q(net310788), .QN(
        n17942) );
  DFF_X1 \REGISTERS_reg[0][29]  ( .D(n3845), .CK(CLK), .Q(net310787), .QN(
        n17941) );
  DFF_X1 \REGISTERS_reg[0][28]  ( .D(n3844), .CK(CLK), .Q(net310786), .QN(
        n17940) );
  DFF_X1 \REGISTERS_reg[0][27]  ( .D(n3843), .CK(CLK), .Q(net310785), .QN(
        n17939) );
  DFF_X1 \REGISTERS_reg[0][26]  ( .D(n3842), .CK(CLK), .Q(net310784), .QN(
        n17938) );
  DFF_X1 \REGISTERS_reg[0][25]  ( .D(n3841), .CK(CLK), .Q(net310783), .QN(
        n17937) );
  DFF_X1 \REGISTERS_reg[0][24]  ( .D(n3840), .CK(CLK), .Q(net310782), .QN(
        n17936) );
  DFF_X1 \REGISTERS_reg[0][23]  ( .D(n3839), .CK(CLK), .Q(net310781), .QN(
        n17967) );
  DFF_X1 \REGISTERS_reg[0][22]  ( .D(n3838), .CK(CLK), .Q(net310780), .QN(
        n17966) );
  DFF_X1 \REGISTERS_reg[0][21]  ( .D(n3837), .CK(CLK), .Q(net310779), .QN(
        n17965) );
  DFF_X1 \REGISTERS_reg[0][20]  ( .D(n3836), .CK(CLK), .Q(net310778), .QN(
        n17964) );
  DFF_X1 \REGISTERS_reg[0][19]  ( .D(n3835), .CK(CLK), .Q(net310777), .QN(
        n17963) );
  DFF_X1 \REGISTERS_reg[0][18]  ( .D(n3834), .CK(CLK), .Q(net310776), .QN(
        n17962) );
  DFF_X1 \REGISTERS_reg[0][17]  ( .D(n3833), .CK(CLK), .Q(net310775), .QN(
        n17961) );
  DFF_X1 \REGISTERS_reg[0][16]  ( .D(n3832), .CK(CLK), .Q(net310774), .QN(
        n17960) );
  DFF_X1 \REGISTERS_reg[0][15]  ( .D(n3831), .CK(CLK), .Q(net310773), .QN(
        n17959) );
  DFF_X1 \REGISTERS_reg[0][14]  ( .D(n3830), .CK(CLK), .Q(net310772), .QN(
        n17958) );
  DFF_X1 \REGISTERS_reg[0][13]  ( .D(n3829), .CK(CLK), .Q(net310771), .QN(
        n17957) );
  DFF_X1 \REGISTERS_reg[0][12]  ( .D(n3828), .CK(CLK), .Q(net310770), .QN(
        n17956) );
  DFF_X1 \REGISTERS_reg[0][11]  ( .D(n3827), .CK(CLK), .Q(net310769), .QN(
        n17955) );
  DFF_X1 \REGISTERS_reg[0][10]  ( .D(n3826), .CK(CLK), .Q(net310768), .QN(
        n17954) );
  DFF_X1 \REGISTERS_reg[0][9]  ( .D(n3825), .CK(CLK), .Q(net310767), .QN(
        n17953) );
  DFF_X1 \REGISTERS_reg[0][8]  ( .D(n3824), .CK(CLK), .Q(net310766), .QN(
        n17952) );
  DFF_X1 \REGISTERS_reg[0][7]  ( .D(n3823), .CK(CLK), .Q(net310765), .QN(
        n17951) );
  DFF_X1 \REGISTERS_reg[0][6]  ( .D(n3822), .CK(CLK), .Q(net310764), .QN(
        n17950) );
  DFF_X1 \REGISTERS_reg[0][5]  ( .D(n3821), .CK(CLK), .Q(net310763), .QN(
        n17949) );
  DFF_X1 \REGISTERS_reg[0][4]  ( .D(n3820), .CK(CLK), .Q(net310762), .QN(
        n17948) );
  DFF_X1 \REGISTERS_reg[0][3]  ( .D(n3819), .CK(CLK), .Q(net310761), .QN(
        n17947) );
  DFF_X1 \REGISTERS_reg[0][2]  ( .D(n3818), .CK(CLK), .Q(net310760), .QN(
        n17946) );
  DFF_X1 \REGISTERS_reg[0][1]  ( .D(n3817), .CK(CLK), .Q(net310759), .QN(
        n17945) );
  DFF_X1 \REGISTERS_reg[0][0]  ( .D(n3816), .CK(CLK), .Q(net310758), .QN(
        n17944) );
  DFF_X1 \REGISTERS_reg[1][31]  ( .D(n3815), .CK(CLK), .Q(net591818), .QN(
        n17726) );
  DFF_X1 \REGISTERS_reg[1][30]  ( .D(n3814), .CK(CLK), .Q(net591817), .QN(
        n17725) );
  DFF_X1 \REGISTERS_reg[1][29]  ( .D(n3813), .CK(CLK), .Q(net591816), .QN(
        n17724) );
  DFF_X1 \REGISTERS_reg[1][28]  ( .D(n3812), .CK(CLK), .Q(net591815), .QN(
        n17723) );
  DFF_X1 \REGISTERS_reg[1][27]  ( .D(n3811), .CK(CLK), .Q(net591814), .QN(
        n17722) );
  DFF_X1 \REGISTERS_reg[1][26]  ( .D(n3810), .CK(CLK), .Q(net591813), .QN(
        n17721) );
  DFF_X1 \REGISTERS_reg[1][25]  ( .D(n3809), .CK(CLK), .Q(net591812), .QN(
        n17720) );
  DFF_X1 \REGISTERS_reg[1][24]  ( .D(n3808), .CK(CLK), .Q(net591811), .QN(
        n17719) );
  DFF_X1 \REGISTERS_reg[1][23]  ( .D(n3807), .CK(CLK), .Q(net591810), .QN(
        n17742) );
  DFF_X1 \REGISTERS_reg[1][22]  ( .D(n3806), .CK(CLK), .Q(net591809), .QN(
        n17741) );
  DFF_X1 \REGISTERS_reg[1][21]  ( .D(n3805), .CK(CLK), .Q(net591808), .QN(
        n17740) );
  DFF_X1 \REGISTERS_reg[1][20]  ( .D(n3804), .CK(CLK), .Q(net591807), .QN(
        n17739) );
  DFF_X1 \REGISTERS_reg[1][19]  ( .D(n3803), .CK(CLK), .Q(net591806), .QN(
        n17738) );
  DFF_X1 \REGISTERS_reg[1][18]  ( .D(n3802), .CK(CLK), .Q(net591805), .QN(
        n17737) );
  DFF_X1 \REGISTERS_reg[1][17]  ( .D(n3801), .CK(CLK), .Q(net591804), .QN(
        n17736) );
  DFF_X1 \REGISTERS_reg[1][16]  ( .D(n3800), .CK(CLK), .Q(net591803), .QN(
        n17735) );
  DFF_X1 \REGISTERS_reg[1][15]  ( .D(n3799), .CK(CLK), .Q(net591802), .QN(
        n17734) );
  DFF_X1 \REGISTERS_reg[1][14]  ( .D(n3798), .CK(CLK), .Q(net591801), .QN(
        n17733) );
  DFF_X1 \REGISTERS_reg[1][13]  ( .D(n3797), .CK(CLK), .Q(net591800), .QN(
        n17732) );
  DFF_X1 \REGISTERS_reg[1][12]  ( .D(n3796), .CK(CLK), .Q(net591799), .QN(
        n17731) );
  DFF_X1 \REGISTERS_reg[1][11]  ( .D(n3795), .CK(CLK), .Q(net591798), .QN(
        n17730) );
  DFF_X1 \REGISTERS_reg[1][10]  ( .D(n3794), .CK(CLK), .Q(net591797), .QN(
        n17729) );
  DFF_X1 \REGISTERS_reg[1][9]  ( .D(n3793), .CK(CLK), .Q(net591796), .QN(
        n17728) );
  DFF_X1 \REGISTERS_reg[1][8]  ( .D(n3792), .CK(CLK), .Q(net591795), .QN(
        n17727) );
  DFF_X1 \REGISTERS_reg[1][7]  ( .D(n3791), .CK(CLK), .Q(net591794), .QN(
        n17718) );
  DFF_X1 \REGISTERS_reg[1][6]  ( .D(n3790), .CK(CLK), .Q(net591793), .QN(
        n17717) );
  DFF_X1 \REGISTERS_reg[1][5]  ( .D(n3789), .CK(CLK), .Q(net591792), .QN(
        n17716) );
  DFF_X1 \REGISTERS_reg[1][4]  ( .D(n3788), .CK(CLK), .Q(net591791), .QN(
        n17714) );
  DFF_X1 \REGISTERS_reg[1][3]  ( .D(n3787), .CK(CLK), .Q(net591790), .QN(
        n17713) );
  DFF_X1 \REGISTERS_reg[1][2]  ( .D(n3786), .CK(CLK), .Q(net591789), .QN(
        n17712) );
  DFF_X1 \REGISTERS_reg[1][1]  ( .D(n3785), .CK(CLK), .Q(net591788), .QN(
        n17711) );
  DFF_X1 \REGISTERS_reg[1][0]  ( .D(n3784), .CK(CLK), .Q(net591787), .QN(
        n17715) );
  DFF_X1 \REGISTERS_reg[2][31]  ( .D(n3783), .CK(CLK), .QN(n17462) );
  DFF_X1 \REGISTERS_reg[2][30]  ( .D(n3782), .CK(CLK), .QN(n17461) );
  DFF_X1 \REGISTERS_reg[2][29]  ( .D(n3781), .CK(CLK), .QN(n17460) );
  DFF_X1 \REGISTERS_reg[2][28]  ( .D(n3780), .CK(CLK), .QN(n17459) );
  DFF_X1 \REGISTERS_reg[2][27]  ( .D(n3779), .CK(CLK), .QN(n17458) );
  DFF_X1 \REGISTERS_reg[2][26]  ( .D(n3778), .CK(CLK), .QN(n17457) );
  DFF_X1 \REGISTERS_reg[2][25]  ( .D(n3777), .CK(CLK), .QN(n17456) );
  DFF_X1 \REGISTERS_reg[2][24]  ( .D(n3776), .CK(CLK), .QN(n17455) );
  DFF_X1 \REGISTERS_reg[2][23]  ( .D(n3775), .CK(CLK), .QN(n17486) );
  DFF_X1 \REGISTERS_reg[2][22]  ( .D(n3774), .CK(CLK), .QN(n17485) );
  DFF_X1 \REGISTERS_reg[2][21]  ( .D(n3773), .CK(CLK), .QN(n17484) );
  DFF_X1 \REGISTERS_reg[2][20]  ( .D(n3772), .CK(CLK), .QN(n17483) );
  DFF_X1 \REGISTERS_reg[2][19]  ( .D(n3771), .CK(CLK), .QN(n17482) );
  DFF_X1 \REGISTERS_reg[2][18]  ( .D(n3770), .CK(CLK), .QN(n17481) );
  DFF_X1 \REGISTERS_reg[2][17]  ( .D(n3769), .CK(CLK), .QN(n17480) );
  DFF_X1 \REGISTERS_reg[2][16]  ( .D(n3768), .CK(CLK), .QN(n17479) );
  DFF_X1 \REGISTERS_reg[2][15]  ( .D(n3767), .CK(CLK), .QN(n17478) );
  DFF_X1 \REGISTERS_reg[2][14]  ( .D(n3766), .CK(CLK), .QN(n17477) );
  DFF_X1 \REGISTERS_reg[2][13]  ( .D(n3765), .CK(CLK), .QN(n17476) );
  DFF_X1 \REGISTERS_reg[2][12]  ( .D(n3764), .CK(CLK), .QN(n17475) );
  DFF_X1 \REGISTERS_reg[2][11]  ( .D(n3763), .CK(CLK), .QN(n17474) );
  DFF_X1 \REGISTERS_reg[2][10]  ( .D(n3762), .CK(CLK), .QN(n17473) );
  DFF_X1 \REGISTERS_reg[2][9]  ( .D(n3761), .CK(CLK), .QN(n17472) );
  DFF_X1 \REGISTERS_reg[2][8]  ( .D(n3760), .CK(CLK), .QN(n17471) );
  DFF_X1 \REGISTERS_reg[2][7]  ( .D(n3759), .CK(CLK), .QN(n17470) );
  DFF_X1 \REGISTERS_reg[2][6]  ( .D(n3758), .CK(CLK), .QN(n17469) );
  DFF_X1 \REGISTERS_reg[2][5]  ( .D(n3757), .CK(CLK), .QN(n17468) );
  DFF_X1 \REGISTERS_reg[2][4]  ( .D(n3756), .CK(CLK), .QN(n17466) );
  DFF_X1 \REGISTERS_reg[2][3]  ( .D(n3755), .CK(CLK), .QN(n17465) );
  DFF_X1 \REGISTERS_reg[2][2]  ( .D(n3754), .CK(CLK), .QN(n17464) );
  DFF_X1 \REGISTERS_reg[2][1]  ( .D(n3753), .CK(CLK), .QN(n17467) );
  DFF_X1 \REGISTERS_reg[2][0]  ( .D(n3752), .CK(CLK), .QN(n17463) );
  DFF_X1 \REGISTERS_reg[3][31]  ( .D(n3751), .CK(CLK), .Q(net423365), .QN(
        n17975) );
  DFF_X1 \REGISTERS_reg[3][30]  ( .D(n3750), .CK(CLK), .Q(net423364), .QN(
        n17974) );
  DFF_X1 \REGISTERS_reg[3][29]  ( .D(n3749), .CK(CLK), .Q(net423363), .QN(
        n17973) );
  DFF_X1 \REGISTERS_reg[3][28]  ( .D(n3748), .CK(CLK), .Q(net423362), .QN(
        n17972) );
  DFF_X1 \REGISTERS_reg[3][27]  ( .D(n3747), .CK(CLK), .Q(net423361), .QN(
        n17971) );
  DFF_X1 \REGISTERS_reg[3][26]  ( .D(n3746), .CK(CLK), .Q(net423360), .QN(
        n17970) );
  DFF_X1 \REGISTERS_reg[3][25]  ( .D(n3745), .CK(CLK), .Q(net423359), .QN(
        n17969) );
  DFF_X1 \REGISTERS_reg[3][24]  ( .D(n3744), .CK(CLK), .Q(net423358), .QN(
        n17968) );
  DFF_X1 \REGISTERS_reg[3][23]  ( .D(n3743), .CK(CLK), .Q(net423357), .QN(
        n17999) );
  DFF_X1 \REGISTERS_reg[3][22]  ( .D(n3742), .CK(CLK), .Q(net423356), .QN(
        n17998) );
  DFF_X1 \REGISTERS_reg[3][21]  ( .D(n3741), .CK(CLK), .Q(net423355), .QN(
        n17997) );
  DFF_X1 \REGISTERS_reg[3][20]  ( .D(n3740), .CK(CLK), .Q(net423354), .QN(
        n17996) );
  DFF_X1 \REGISTERS_reg[3][19]  ( .D(n3739), .CK(CLK), .Q(net423353), .QN(
        n17995) );
  DFF_X1 \REGISTERS_reg[3][18]  ( .D(n3738), .CK(CLK), .Q(net423352), .QN(
        n17994) );
  DFF_X1 \REGISTERS_reg[3][17]  ( .D(n3737), .CK(CLK), .Q(net423351), .QN(
        n17993) );
  DFF_X1 \REGISTERS_reg[3][16]  ( .D(n3736), .CK(CLK), .Q(net423350), .QN(
        n17992) );
  DFF_X1 \REGISTERS_reg[3][15]  ( .D(n3735), .CK(CLK), .Q(net423349), .QN(
        n17991) );
  DFF_X1 \REGISTERS_reg[3][14]  ( .D(n3734), .CK(CLK), .Q(net423348), .QN(
        n17990) );
  DFF_X1 \REGISTERS_reg[3][13]  ( .D(n3733), .CK(CLK), .Q(net423347), .QN(
        n17989) );
  DFF_X1 \REGISTERS_reg[3][12]  ( .D(n3732), .CK(CLK), .Q(net423346), .QN(
        n17988) );
  DFF_X1 \REGISTERS_reg[3][11]  ( .D(n3731), .CK(CLK), .Q(net423345), .QN(
        n17987) );
  DFF_X1 \REGISTERS_reg[3][10]  ( .D(n3730), .CK(CLK), .Q(net423344), .QN(
        n17986) );
  DFF_X1 \REGISTERS_reg[3][9]  ( .D(n3729), .CK(CLK), .Q(net423343), .QN(
        n17985) );
  DFF_X1 \REGISTERS_reg[3][8]  ( .D(n3728), .CK(CLK), .Q(net423342), .QN(
        n17984) );
  DFF_X1 \REGISTERS_reg[3][7]  ( .D(n3727), .CK(CLK), .Q(net423341), .QN(
        n17983) );
  DFF_X1 \REGISTERS_reg[3][6]  ( .D(n3726), .CK(CLK), .Q(net423340), .QN(
        n17982) );
  DFF_X1 \REGISTERS_reg[3][5]  ( .D(n3725), .CK(CLK), .Q(net423339), .QN(
        n17981) );
  DFF_X1 \REGISTERS_reg[3][4]  ( .D(n3724), .CK(CLK), .Q(net423338), .QN(
        n17978) );
  DFF_X1 \REGISTERS_reg[3][3]  ( .D(n3723), .CK(CLK), .Q(net423337), .QN(
        n17977) );
  DFF_X1 \REGISTERS_reg[3][2]  ( .D(n3722), .CK(CLK), .Q(net423336), .QN(
        n17976) );
  DFF_X1 \REGISTERS_reg[3][1]  ( .D(n3721), .CK(CLK), .Q(net423335), .QN(
        n17980) );
  DFF_X1 \REGISTERS_reg[3][0]  ( .D(n3720), .CK(CLK), .Q(net423334), .QN(
        n17979) );
  DFF_X1 \REGISTERS_reg[4][31]  ( .D(n3719), .CK(CLK), .Q(net591754), .QN(
        n18261) );
  DFF_X1 \REGISTERS_reg[4][30]  ( .D(n3718), .CK(CLK), .Q(net591753), .QN(
        n18260) );
  DFF_X1 \REGISTERS_reg[4][29]  ( .D(n3717), .CK(CLK), .Q(net591752), .QN(
        n18259) );
  DFF_X1 \REGISTERS_reg[4][28]  ( .D(n3716), .CK(CLK), .Q(net591751), .QN(
        n18258) );
  DFF_X1 \REGISTERS_reg[4][27]  ( .D(n3715), .CK(CLK), .Q(net591750), .QN(
        n18257) );
  DFF_X1 \REGISTERS_reg[4][26]  ( .D(n3714), .CK(CLK), .Q(net591749), .QN(
        n18256) );
  DFF_X1 \REGISTERS_reg[4][25]  ( .D(n3713), .CK(CLK), .Q(net591748), .QN(
        n18255) );
  DFF_X1 \REGISTERS_reg[4][24]  ( .D(n3712), .CK(CLK), .Q(net591747), .QN(
        n18254) );
  DFF_X1 \REGISTERS_reg[4][23]  ( .D(n3711), .CK(CLK), .Q(net591746), .QN(
        n18285) );
  DFF_X1 \REGISTERS_reg[4][22]  ( .D(n3710), .CK(CLK), .Q(net591745), .QN(
        n18284) );
  DFF_X1 \REGISTERS_reg[4][21]  ( .D(n3709), .CK(CLK), .Q(net591744), .QN(
        n18283) );
  DFF_X1 \REGISTERS_reg[4][20]  ( .D(n3708), .CK(CLK), .Q(net591743), .QN(
        n18282) );
  DFF_X1 \REGISTERS_reg[4][19]  ( .D(n3707), .CK(CLK), .Q(net591742), .QN(
        n18281) );
  DFF_X1 \REGISTERS_reg[4][18]  ( .D(n3706), .CK(CLK), .Q(net591741), .QN(
        n18280) );
  DFF_X1 \REGISTERS_reg[4][17]  ( .D(n3705), .CK(CLK), .Q(net591740), .QN(
        n18279) );
  DFF_X1 \REGISTERS_reg[4][16]  ( .D(n3704), .CK(CLK), .Q(net591739), .QN(
        n18278) );
  DFF_X1 \REGISTERS_reg[4][15]  ( .D(n3703), .CK(CLK), .Q(net591738), .QN(
        n18277) );
  DFF_X1 \REGISTERS_reg[4][14]  ( .D(n3702), .CK(CLK), .Q(net591737), .QN(
        n18276) );
  DFF_X1 \REGISTERS_reg[4][13]  ( .D(n3701), .CK(CLK), .Q(net591736), .QN(
        n18275) );
  DFF_X1 \REGISTERS_reg[4][12]  ( .D(n3700), .CK(CLK), .Q(net591735), .QN(
        n18274) );
  DFF_X1 \REGISTERS_reg[4][11]  ( .D(n3699), .CK(CLK), .Q(net591734), .QN(
        n18273) );
  DFF_X1 \REGISTERS_reg[4][10]  ( .D(n3698), .CK(CLK), .Q(net591733), .QN(
        n18272) );
  DFF_X1 \REGISTERS_reg[4][9]  ( .D(n3697), .CK(CLK), .Q(net591732), .QN(
        n18271) );
  DFF_X1 \REGISTERS_reg[4][8]  ( .D(n3696), .CK(CLK), .Q(net591731), .QN(
        n18270) );
  DFF_X1 \REGISTERS_reg[4][7]  ( .D(n3695), .CK(CLK), .Q(net591730), .QN(
        n18269) );
  DFF_X1 \REGISTERS_reg[4][6]  ( .D(n3694), .CK(CLK), .Q(net591729), .QN(
        n18268) );
  DFF_X1 \REGISTERS_reg[4][5]  ( .D(n3693), .CK(CLK), .Q(net591728), .QN(
        n18267) );
  DFF_X1 \REGISTERS_reg[4][4]  ( .D(n3692), .CK(CLK), .Q(net591727), .QN(
        n18265) );
  DFF_X1 \REGISTERS_reg[4][3]  ( .D(n3691), .CK(CLK), .Q(net591726), .QN(
        n18264) );
  DFF_X1 \REGISTERS_reg[4][2]  ( .D(n3690), .CK(CLK), .Q(net591725), .QN(
        n18266) );
  DFF_X1 \REGISTERS_reg[4][1]  ( .D(n3689), .CK(CLK), .Q(net591724), .QN(
        n18263) );
  DFF_X1 \REGISTERS_reg[4][0]  ( .D(n3688), .CK(CLK), .Q(net591723), .QN(
        n18262) );
  DFF_X1 \REGISTERS_reg[5][31]  ( .D(n3687), .CK(CLK), .Q(net367142), .QN(
        n18015) );
  DFF_X1 \REGISTERS_reg[5][30]  ( .D(n3686), .CK(CLK), .Q(net367141), .QN(
        n18014) );
  DFF_X1 \REGISTERS_reg[5][29]  ( .D(n3685), .CK(CLK), .Q(net367140), .QN(
        n18013) );
  DFF_X1 \REGISTERS_reg[5][28]  ( .D(n3684), .CK(CLK), .Q(net367139), .QN(
        n18012) );
  DFF_X1 \REGISTERS_reg[5][27]  ( .D(n3683), .CK(CLK), .Q(net367138), .QN(
        n18011) );
  DFF_X1 \REGISTERS_reg[5][26]  ( .D(n3682), .CK(CLK), .Q(net367137), .QN(
        n18010) );
  DFF_X1 \REGISTERS_reg[5][25]  ( .D(n3681), .CK(CLK), .Q(net367136), .QN(
        n18009) );
  DFF_X1 \REGISTERS_reg[5][24]  ( .D(n3680), .CK(CLK), .Q(net367135), .QN(
        n18008) );
  DFF_X1 \REGISTERS_reg[5][23]  ( .D(n3679), .CK(CLK), .Q(net367134), .QN(
        n18063) );
  DFF_X1 \REGISTERS_reg[5][22]  ( .D(n3678), .CK(CLK), .Q(net367133), .QN(
        n18062) );
  DFF_X1 \REGISTERS_reg[5][21]  ( .D(n3677), .CK(CLK), .Q(net367132), .QN(
        n18061) );
  DFF_X1 \REGISTERS_reg[5][20]  ( .D(n3676), .CK(CLK), .Q(net367131), .QN(
        n18060) );
  DFF_X1 \REGISTERS_reg[5][19]  ( .D(n3675), .CK(CLK), .Q(net367130), .QN(
        n18059) );
  DFF_X1 \REGISTERS_reg[5][18]  ( .D(n3674), .CK(CLK), .Q(net367129), .QN(
        n18058) );
  DFF_X1 \REGISTERS_reg[5][17]  ( .D(n3673), .CK(CLK), .Q(net367128), .QN(
        n18057) );
  DFF_X1 \REGISTERS_reg[5][16]  ( .D(n3672), .CK(CLK), .Q(net367127), .QN(
        n18056) );
  DFF_X1 \REGISTERS_reg[5][15]  ( .D(n3671), .CK(CLK), .Q(net367126), .QN(
        n18055) );
  DFF_X1 \REGISTERS_reg[5][14]  ( .D(n3670), .CK(CLK), .Q(net367125), .QN(
        n18054) );
  DFF_X1 \REGISTERS_reg[5][13]  ( .D(n3669), .CK(CLK), .Q(net367124), .QN(
        n18053) );
  DFF_X1 \REGISTERS_reg[5][12]  ( .D(n3668), .CK(CLK), .Q(net367123), .QN(
        n18052) );
  DFF_X1 \REGISTERS_reg[5][11]  ( .D(n3667), .CK(CLK), .Q(net367122), .QN(
        n18051) );
  DFF_X1 \REGISTERS_reg[5][10]  ( .D(n3666), .CK(CLK), .Q(net367121), .QN(
        n18050) );
  DFF_X1 \REGISTERS_reg[5][9]  ( .D(n3665), .CK(CLK), .Q(net367120), .QN(
        n18049) );
  DFF_X1 \REGISTERS_reg[5][8]  ( .D(n3664), .CK(CLK), .Q(net367119), .QN(
        n18048) );
  DFF_X1 \REGISTERS_reg[5][7]  ( .D(n3663), .CK(CLK), .Q(net367118), .QN(
        n18047) );
  DFF_X1 \REGISTERS_reg[5][6]  ( .D(n3662), .CK(CLK), .Q(net367117), .QN(
        n18046) );
  DFF_X1 \REGISTERS_reg[5][5]  ( .D(n3661), .CK(CLK), .Q(net367116), .QN(
        n18045) );
  DFF_X1 \REGISTERS_reg[5][4]  ( .D(n3660), .CK(CLK), .Q(net367115), .QN(
        n18021) );
  DFF_X1 \REGISTERS_reg[5][3]  ( .D(n3659), .CK(CLK), .Q(net367114), .QN(
        n18020) );
  DFF_X1 \REGISTERS_reg[5][2]  ( .D(n3658), .CK(CLK), .Q(net367113), .QN(
        n18044) );
  DFF_X1 \REGISTERS_reg[5][1]  ( .D(n3657), .CK(CLK), .Q(net367112), .QN(
        n18019) );
  DFF_X1 \REGISTERS_reg[5][0]  ( .D(n3656), .CK(CLK), .Q(net367111), .QN(
        n18043) );
  DFF_X1 \REGISTERS_reg[6][31]  ( .D(n3655), .CK(CLK), .QN(n17334) );
  DFF_X1 \REGISTERS_reg[6][30]  ( .D(n3654), .CK(CLK), .QN(n17333) );
  DFF_X1 \REGISTERS_reg[6][29]  ( .D(n3653), .CK(CLK), .QN(n17332) );
  DFF_X1 \REGISTERS_reg[6][28]  ( .D(n3652), .CK(CLK), .QN(n17331) );
  DFF_X1 \REGISTERS_reg[6][27]  ( .D(n3651), .CK(CLK), .QN(n17330) );
  DFF_X1 \REGISTERS_reg[6][26]  ( .D(n3650), .CK(CLK), .QN(n17329) );
  DFF_X1 \REGISTERS_reg[6][25]  ( .D(n3649), .CK(CLK), .QN(n17328) );
  DFF_X1 \REGISTERS_reg[6][24]  ( .D(n3648), .CK(CLK), .QN(n17327) );
  DFF_X1 \REGISTERS_reg[6][23]  ( .D(n3647), .CK(CLK), .QN(n17358) );
  DFF_X1 \REGISTERS_reg[6][22]  ( .D(n3646), .CK(CLK), .QN(n17357) );
  DFF_X1 \REGISTERS_reg[6][21]  ( .D(n3645), .CK(CLK), .QN(n17356) );
  DFF_X1 \REGISTERS_reg[6][20]  ( .D(n3644), .CK(CLK), .QN(n17355) );
  DFF_X1 \REGISTERS_reg[6][19]  ( .D(n3643), .CK(CLK), .QN(n17354) );
  DFF_X1 \REGISTERS_reg[6][18]  ( .D(n3642), .CK(CLK), .QN(n17353) );
  DFF_X1 \REGISTERS_reg[6][17]  ( .D(n3641), .CK(CLK), .QN(n17352) );
  DFF_X1 \REGISTERS_reg[6][16]  ( .D(n3640), .CK(CLK), .QN(n17351) );
  DFF_X1 \REGISTERS_reg[6][15]  ( .D(n3639), .CK(CLK), .QN(n17350) );
  DFF_X1 \REGISTERS_reg[6][14]  ( .D(n3638), .CK(CLK), .QN(n17349) );
  DFF_X1 \REGISTERS_reg[6][13]  ( .D(n3637), .CK(CLK), .QN(n17348) );
  DFF_X1 \REGISTERS_reg[6][12]  ( .D(n3636), .CK(CLK), .QN(n17347) );
  DFF_X1 \REGISTERS_reg[6][11]  ( .D(n3635), .CK(CLK), .QN(n17346) );
  DFF_X1 \REGISTERS_reg[6][10]  ( .D(n3634), .CK(CLK), .QN(n17345) );
  DFF_X1 \REGISTERS_reg[6][9]  ( .D(n3633), .CK(CLK), .QN(n17344) );
  DFF_X1 \REGISTERS_reg[6][8]  ( .D(n3632), .CK(CLK), .QN(n17343) );
  DFF_X1 \REGISTERS_reg[6][7]  ( .D(n3631), .CK(CLK), .QN(n17342) );
  DFF_X1 \REGISTERS_reg[6][6]  ( .D(n3630), .CK(CLK), .QN(n17341) );
  DFF_X1 \REGISTERS_reg[6][5]  ( .D(n3629), .CK(CLK), .QN(n17340) );
  DFF_X1 \REGISTERS_reg[6][4]  ( .D(n3628), .CK(CLK), .QN(n17337) );
  DFF_X1 \REGISTERS_reg[6][3]  ( .D(n3627), .CK(CLK), .QN(n17336) );
  DFF_X1 \REGISTERS_reg[6][2]  ( .D(n3626), .CK(CLK), .QN(n17339) );
  DFF_X1 \REGISTERS_reg[6][1]  ( .D(n3625), .CK(CLK), .QN(n17338) );
  DFF_X1 \REGISTERS_reg[6][0]  ( .D(n3624), .CK(CLK), .QN(n17335) );
  DFF_X1 \REGISTERS_reg[7][31]  ( .D(n3623), .CK(CLK), .Q(net535563), .QN(
        n17814) );
  DFF_X1 \REGISTERS_reg[7][30]  ( .D(n3622), .CK(CLK), .Q(net535562), .QN(
        n17813) );
  DFF_X1 \REGISTERS_reg[7][29]  ( .D(n3621), .CK(CLK), .Q(net535561), .QN(
        n17812) );
  DFF_X1 \REGISTERS_reg[7][28]  ( .D(n3620), .CK(CLK), .Q(net535560), .QN(
        n17811) );
  DFF_X1 \REGISTERS_reg[7][27]  ( .D(n3619), .CK(CLK), .Q(net535559), .QN(
        n17810) );
  DFF_X1 \REGISTERS_reg[7][26]  ( .D(n3618), .CK(CLK), .Q(net535558), .QN(
        n17809) );
  DFF_X1 \REGISTERS_reg[7][25]  ( .D(n3617), .CK(CLK), .Q(net535557), .QN(
        n17808) );
  DFF_X1 \REGISTERS_reg[7][24]  ( .D(n3616), .CK(CLK), .Q(net535556), .QN(
        n17807) );
  DFF_X1 \REGISTERS_reg[7][23]  ( .D(n3615), .CK(CLK), .Q(net535555), .QN(
        n17838) );
  DFF_X1 \REGISTERS_reg[7][22]  ( .D(n3614), .CK(CLK), .Q(net535554), .QN(
        n17837) );
  DFF_X1 \REGISTERS_reg[7][21]  ( .D(n3613), .CK(CLK), .Q(net535553), .QN(
        n17836) );
  DFF_X1 \REGISTERS_reg[7][20]  ( .D(n3612), .CK(CLK), .Q(net535552), .QN(
        n17835) );
  DFF_X1 \REGISTERS_reg[7][19]  ( .D(n3611), .CK(CLK), .Q(net535551), .QN(
        n17834) );
  DFF_X1 \REGISTERS_reg[7][18]  ( .D(n3610), .CK(CLK), .Q(net535550), .QN(
        n17833) );
  DFF_X1 \REGISTERS_reg[7][17]  ( .D(n3609), .CK(CLK), .Q(net535549), .QN(
        n17832) );
  DFF_X1 \REGISTERS_reg[7][16]  ( .D(n3608), .CK(CLK), .Q(net535548), .QN(
        n17831) );
  DFF_X1 \REGISTERS_reg[7][15]  ( .D(n3607), .CK(CLK), .Q(net535547), .QN(
        n17830) );
  DFF_X1 \REGISTERS_reg[7][14]  ( .D(n3606), .CK(CLK), .Q(net535546), .QN(
        n17829) );
  DFF_X1 \REGISTERS_reg[7][13]  ( .D(n3605), .CK(CLK), .Q(net535545), .QN(
        n17828) );
  DFF_X1 \REGISTERS_reg[7][12]  ( .D(n3604), .CK(CLK), .Q(net535544), .QN(
        n17827) );
  DFF_X1 \REGISTERS_reg[7][11]  ( .D(n3603), .CK(CLK), .Q(net535543), .QN(
        n17826) );
  DFF_X1 \REGISTERS_reg[7][10]  ( .D(n3602), .CK(CLK), .Q(net535542), .QN(
        n17825) );
  DFF_X1 \REGISTERS_reg[7][9]  ( .D(n3601), .CK(CLK), .Q(net535541), .QN(
        n17824) );
  DFF_X1 \REGISTERS_reg[7][8]  ( .D(n3600), .CK(CLK), .Q(net535540), .QN(
        n17823) );
  DFF_X1 \REGISTERS_reg[7][7]  ( .D(n3599), .CK(CLK), .Q(net535539), .QN(
        n17822) );
  DFF_X1 \REGISTERS_reg[7][6]  ( .D(n3598), .CK(CLK), .Q(net535538), .QN(
        n17821) );
  DFF_X1 \REGISTERS_reg[7][5]  ( .D(n3597), .CK(CLK), .Q(net535537), .QN(
        n17820) );
  DFF_X1 \REGISTERS_reg[7][4]  ( .D(n3596), .CK(CLK), .Q(net535536), .QN(
        n17816) );
  DFF_X1 \REGISTERS_reg[7][3]  ( .D(n3595), .CK(CLK), .Q(net535535), .QN(
        n17815) );
  DFF_X1 \REGISTERS_reg[7][2]  ( .D(n3594), .CK(CLK), .Q(net535534), .QN(
        n17819) );
  DFF_X1 \REGISTERS_reg[7][1]  ( .D(n3593), .CK(CLK), .Q(net535533), .QN(
        n17818) );
  DFF_X1 \REGISTERS_reg[7][0]  ( .D(n3592), .CK(CLK), .Q(net535532), .QN(
        n17817) );
  DFF_X1 \REGISTERS_reg[8][31]  ( .D(n3591), .CK(CLK), .Q(net535531), .QN(
        n17686) );
  DFF_X1 \REGISTERS_reg[8][30]  ( .D(n3590), .CK(CLK), .Q(net535530), .QN(
        n17685) );
  DFF_X1 \REGISTERS_reg[8][29]  ( .D(n3589), .CK(CLK), .Q(net535529), .QN(
        n17684) );
  DFF_X1 \REGISTERS_reg[8][28]  ( .D(n3588), .CK(CLK), .Q(net535528), .QN(
        n17683) );
  DFF_X1 \REGISTERS_reg[8][27]  ( .D(n3587), .CK(CLK), .Q(net535527), .QN(
        n17682) );
  DFF_X1 \REGISTERS_reg[8][26]  ( .D(n3586), .CK(CLK), .Q(net535526), .QN(
        n17681) );
  DFF_X1 \REGISTERS_reg[8][25]  ( .D(n3585), .CK(CLK), .Q(net535525), .QN(
        n17680) );
  DFF_X1 \REGISTERS_reg[8][24]  ( .D(n3584), .CK(CLK), .Q(net535524), .QN(
        n17679) );
  DFF_X1 \REGISTERS_reg[8][23]  ( .D(n3583), .CK(CLK), .Q(net535523), .QN(
        n17710) );
  DFF_X1 \REGISTERS_reg[8][22]  ( .D(n3582), .CK(CLK), .Q(net535522), .QN(
        n17709) );
  DFF_X1 \REGISTERS_reg[8][21]  ( .D(n3581), .CK(CLK), .Q(net535521), .QN(
        n17708) );
  DFF_X1 \REGISTERS_reg[8][20]  ( .D(n3580), .CK(CLK), .Q(net535520), .QN(
        n17707) );
  DFF_X1 \REGISTERS_reg[8][19]  ( .D(n3579), .CK(CLK), .Q(net535519), .QN(
        n17706) );
  DFF_X1 \REGISTERS_reg[8][18]  ( .D(n3578), .CK(CLK), .Q(net535518), .QN(
        n17705) );
  DFF_X1 \REGISTERS_reg[8][17]  ( .D(n3577), .CK(CLK), .Q(net535517), .QN(
        n17704) );
  DFF_X1 \REGISTERS_reg[8][16]  ( .D(n3576), .CK(CLK), .Q(net535516), .QN(
        n17703) );
  DFF_X1 \REGISTERS_reg[8][15]  ( .D(n3575), .CK(CLK), .Q(net535515), .QN(
        n17702) );
  DFF_X1 \REGISTERS_reg[8][14]  ( .D(n3574), .CK(CLK), .Q(net535514), .QN(
        n17701) );
  DFF_X1 \REGISTERS_reg[8][13]  ( .D(n3573), .CK(CLK), .Q(net535513), .QN(
        n17700) );
  DFF_X1 \REGISTERS_reg[8][12]  ( .D(n3572), .CK(CLK), .Q(net535512), .QN(
        n17699) );
  DFF_X1 \REGISTERS_reg[8][11]  ( .D(n3571), .CK(CLK), .Q(net535511), .QN(
        n17698) );
  DFF_X1 \REGISTERS_reg[8][10]  ( .D(n3570), .CK(CLK), .Q(net535510), .QN(
        n17697) );
  DFF_X1 \REGISTERS_reg[8][9]  ( .D(n3569), .CK(CLK), .Q(net535509), .QN(
        n17696) );
  DFF_X1 \REGISTERS_reg[8][8]  ( .D(n3568), .CK(CLK), .Q(net535508), .QN(
        n17695) );
  DFF_X1 \REGISTERS_reg[8][7]  ( .D(n3567), .CK(CLK), .Q(net535507), .QN(
        n17694) );
  DFF_X1 \REGISTERS_reg[8][6]  ( .D(n3566), .CK(CLK), .Q(net535506), .QN(
        n17693) );
  DFF_X1 \REGISTERS_reg[8][5]  ( .D(n3565), .CK(CLK), .Q(net535505), .QN(
        n17692) );
  DFF_X1 \REGISTERS_reg[8][4]  ( .D(n3564), .CK(CLK), .Q(net535504), .QN(
        n17690) );
  DFF_X1 \REGISTERS_reg[8][3]  ( .D(n3563), .CK(CLK), .Q(net535503), .QN(
        n17691) );
  DFF_X1 \REGISTERS_reg[8][2]  ( .D(n3562), .CK(CLK), .Q(net535502), .QN(
        n17689) );
  DFF_X1 \REGISTERS_reg[8][1]  ( .D(n3561), .CK(CLK), .Q(net535501), .QN(
        n17688) );
  DFF_X1 \REGISTERS_reg[8][0]  ( .D(n3560), .CK(CLK), .Q(net535500), .QN(
        n17687) );
  DFF_X1 \REGISTERS_reg[9][31]  ( .D(n3559), .CK(CLK), .QN(n17398) );
  DFF_X1 \REGISTERS_reg[9][30]  ( .D(n3558), .CK(CLK), .QN(n17397) );
  DFF_X1 \REGISTERS_reg[9][29]  ( .D(n3557), .CK(CLK), .QN(n17396) );
  DFF_X1 \REGISTERS_reg[9][28]  ( .D(n3556), .CK(CLK), .QN(n17395) );
  DFF_X1 \REGISTERS_reg[9][27]  ( .D(n3555), .CK(CLK), .QN(n17394) );
  DFF_X1 \REGISTERS_reg[9][26]  ( .D(n3554), .CK(CLK), .QN(n17393) );
  DFF_X1 \REGISTERS_reg[9][25]  ( .D(n3553), .CK(CLK), .QN(n17392) );
  DFF_X1 \REGISTERS_reg[9][24]  ( .D(n3552), .CK(CLK), .QN(n17391) );
  DFF_X1 \REGISTERS_reg[9][23]  ( .D(n3551), .CK(CLK), .QN(n17422) );
  DFF_X1 \REGISTERS_reg[9][22]  ( .D(n3550), .CK(CLK), .QN(n17421) );
  DFF_X1 \REGISTERS_reg[9][21]  ( .D(n3549), .CK(CLK), .QN(n17420) );
  DFF_X1 \REGISTERS_reg[9][20]  ( .D(n3548), .CK(CLK), .QN(n17419) );
  DFF_X1 \REGISTERS_reg[9][19]  ( .D(n3547), .CK(CLK), .QN(n17418) );
  DFF_X1 \REGISTERS_reg[9][18]  ( .D(n3546), .CK(CLK), .QN(n17417) );
  DFF_X1 \REGISTERS_reg[9][17]  ( .D(n3545), .CK(CLK), .QN(n17416) );
  DFF_X1 \REGISTERS_reg[9][16]  ( .D(n3544), .CK(CLK), .QN(n17415) );
  DFF_X1 \REGISTERS_reg[9][15]  ( .D(n3543), .CK(CLK), .QN(n17414) );
  DFF_X1 \REGISTERS_reg[9][14]  ( .D(n3542), .CK(CLK), .QN(n17413) );
  DFF_X1 \REGISTERS_reg[9][13]  ( .D(n3541), .CK(CLK), .QN(n17412) );
  DFF_X1 \REGISTERS_reg[9][12]  ( .D(n3540), .CK(CLK), .QN(n17411) );
  DFF_X1 \REGISTERS_reg[9][11]  ( .D(n3539), .CK(CLK), .QN(n17410) );
  DFF_X1 \REGISTERS_reg[9][10]  ( .D(n3538), .CK(CLK), .QN(n17409) );
  DFF_X1 \REGISTERS_reg[9][9]  ( .D(n3537), .CK(CLK), .QN(n17408) );
  DFF_X1 \REGISTERS_reg[9][8]  ( .D(n3536), .CK(CLK), .QN(n17407) );
  DFF_X1 \REGISTERS_reg[9][7]  ( .D(n3535), .CK(CLK), .QN(n17406) );
  DFF_X1 \REGISTERS_reg[9][6]  ( .D(n3534), .CK(CLK), .QN(n17405) );
  DFF_X1 \REGISTERS_reg[9][5]  ( .D(n3533), .CK(CLK), .QN(n17404) );
  DFF_X1 \REGISTERS_reg[9][4]  ( .D(n3532), .CK(CLK), .QN(n17401) );
  DFF_X1 \REGISTERS_reg[9][3]  ( .D(n3531), .CK(CLK), .QN(n17403) );
  DFF_X1 \REGISTERS_reg[9][2]  ( .D(n3530), .CK(CLK), .QN(n17400) );
  DFF_X1 \REGISTERS_reg[9][1]  ( .D(n3529), .CK(CLK), .QN(n17399) );
  DFF_X1 \REGISTERS_reg[9][0]  ( .D(n3528), .CK(CLK), .QN(n17402) );
  DFF_X1 \REGISTERS_reg[10][31]  ( .D(n3527), .CK(CLK), .QN(n17534) );
  DFF_X1 \REGISTERS_reg[10][30]  ( .D(n3526), .CK(CLK), .QN(n17533) );
  DFF_X1 \REGISTERS_reg[10][29]  ( .D(n3525), .CK(CLK), .QN(n17532) );
  DFF_X1 \REGISTERS_reg[10][28]  ( .D(n3524), .CK(CLK), .QN(n17531) );
  DFF_X1 \REGISTERS_reg[10][27]  ( .D(n3523), .CK(CLK), .QN(n17530) );
  DFF_X1 \REGISTERS_reg[10][26]  ( .D(n3522), .CK(CLK), .QN(n17529) );
  DFF_X1 \REGISTERS_reg[10][25]  ( .D(n3521), .CK(CLK), .QN(n17528) );
  DFF_X1 \REGISTERS_reg[10][24]  ( .D(n3520), .CK(CLK), .QN(n17527) );
  DFF_X1 \REGISTERS_reg[10][23]  ( .D(n3519), .CK(CLK), .QN(n17582) );
  DFF_X1 \REGISTERS_reg[10][22]  ( .D(n3518), .CK(CLK), .QN(n17581) );
  DFF_X1 \REGISTERS_reg[10][21]  ( .D(n3517), .CK(CLK), .QN(n17580) );
  DFF_X1 \REGISTERS_reg[10][20]  ( .D(n3516), .CK(CLK), .QN(n17579) );
  DFF_X1 \REGISTERS_reg[10][19]  ( .D(n3515), .CK(CLK), .QN(n17578) );
  DFF_X1 \REGISTERS_reg[10][18]  ( .D(n3514), .CK(CLK), .QN(n17577) );
  DFF_X1 \REGISTERS_reg[10][17]  ( .D(n3513), .CK(CLK), .QN(n17576) );
  DFF_X1 \REGISTERS_reg[10][16]  ( .D(n3512), .CK(CLK), .QN(n17575) );
  DFF_X1 \REGISTERS_reg[10][15]  ( .D(n3511), .CK(CLK), .QN(n17574) );
  DFF_X1 \REGISTERS_reg[10][14]  ( .D(n3510), .CK(CLK), .QN(n17573) );
  DFF_X1 \REGISTERS_reg[10][13]  ( .D(n3509), .CK(CLK), .QN(n17572) );
  DFF_X1 \REGISTERS_reg[10][12]  ( .D(n3508), .CK(CLK), .QN(n17571) );
  DFF_X1 \REGISTERS_reg[10][11]  ( .D(n3507), .CK(CLK), .QN(n17570) );
  DFF_X1 \REGISTERS_reg[10][10]  ( .D(n3506), .CK(CLK), .QN(n17569) );
  DFF_X1 \REGISTERS_reg[10][9]  ( .D(n3505), .CK(CLK), .QN(n17568) );
  DFF_X1 \REGISTERS_reg[10][8]  ( .D(n3504), .CK(CLK), .QN(n17567) );
  DFF_X1 \REGISTERS_reg[10][7]  ( .D(n3503), .CK(CLK), .QN(n17566) );
  DFF_X1 \REGISTERS_reg[10][6]  ( .D(n3502), .CK(CLK), .QN(n17565) );
  DFF_X1 \REGISTERS_reg[10][5]  ( .D(n3501), .CK(CLK), .QN(n17564) );
  DFF_X1 \REGISTERS_reg[10][4]  ( .D(n3500), .CK(CLK), .QN(n17539) );
  DFF_X1 \REGISTERS_reg[10][3]  ( .D(n3499), .CK(CLK), .QN(n17563) );
  DFF_X1 \REGISTERS_reg[10][2]  ( .D(n3498), .CK(CLK), .QN(n17538) );
  DFF_X1 \REGISTERS_reg[10][1]  ( .D(n3497), .CK(CLK), .QN(n17562) );
  DFF_X1 \REGISTERS_reg[10][0]  ( .D(n3496), .CK(CLK), .QN(n17537) );
  DFF_X1 \REGISTERS_reg[11][31]  ( .D(n3495), .CK(CLK), .Q(net479441), .QN(
        n18079) );
  DFF_X1 \REGISTERS_reg[11][30]  ( .D(n3494), .CK(CLK), .Q(net479440), .QN(
        n18078) );
  DFF_X1 \REGISTERS_reg[11][29]  ( .D(n3493), .CK(CLK), .Q(net479439), .QN(
        n18077) );
  DFF_X1 \REGISTERS_reg[11][28]  ( .D(n3492), .CK(CLK), .Q(net479438), .QN(
        n18076) );
  DFF_X1 \REGISTERS_reg[11][27]  ( .D(n3491), .CK(CLK), .Q(net479437), .QN(
        n18075) );
  DFF_X1 \REGISTERS_reg[11][26]  ( .D(n3490), .CK(CLK), .Q(net479436), .QN(
        n18074) );
  DFF_X1 \REGISTERS_reg[11][25]  ( .D(n3489), .CK(CLK), .Q(net479435), .QN(
        n18073) );
  DFF_X1 \REGISTERS_reg[11][24]  ( .D(n3488), .CK(CLK), .Q(net479434), .QN(
        n18072) );
  DFF_X1 \REGISTERS_reg[11][23]  ( .D(n3487), .CK(CLK), .Q(net479433), .QN(
        n18127) );
  DFF_X1 \REGISTERS_reg[11][22]  ( .D(n3486), .CK(CLK), .Q(net479432), .QN(
        n18126) );
  DFF_X1 \REGISTERS_reg[11][21]  ( .D(n3485), .CK(CLK), .Q(net479431), .QN(
        n18125) );
  DFF_X1 \REGISTERS_reg[11][20]  ( .D(n3484), .CK(CLK), .Q(net479430), .QN(
        n18124) );
  DFF_X1 \REGISTERS_reg[11][19]  ( .D(n3483), .CK(CLK), .Q(net479429), .QN(
        n18123) );
  DFF_X1 \REGISTERS_reg[11][18]  ( .D(n3482), .CK(CLK), .Q(net479428), .QN(
        n18122) );
  DFF_X1 \REGISTERS_reg[11][17]  ( .D(n3481), .CK(CLK), .Q(net479427), .QN(
        n18121) );
  DFF_X1 \REGISTERS_reg[11][16]  ( .D(n3480), .CK(CLK), .Q(net479426), .QN(
        n18120) );
  DFF_X1 \REGISTERS_reg[11][15]  ( .D(n3479), .CK(CLK), .Q(net479425), .QN(
        n18119) );
  DFF_X1 \REGISTERS_reg[11][14]  ( .D(n3478), .CK(CLK), .Q(net479424), .QN(
        n18118) );
  DFF_X1 \REGISTERS_reg[11][13]  ( .D(n3477), .CK(CLK), .Q(net479423), .QN(
        n18117) );
  DFF_X1 \REGISTERS_reg[11][12]  ( .D(n3476), .CK(CLK), .Q(net479422), .QN(
        n18116) );
  DFF_X1 \REGISTERS_reg[11][11]  ( .D(n3475), .CK(CLK), .Q(net479421), .QN(
        n18115) );
  DFF_X1 \REGISTERS_reg[11][10]  ( .D(n3474), .CK(CLK), .Q(net479420), .QN(
        n18114) );
  DFF_X1 \REGISTERS_reg[11][9]  ( .D(n3473), .CK(CLK), .Q(net479419), .QN(
        n18113) );
  DFF_X1 \REGISTERS_reg[11][8]  ( .D(n3472), .CK(CLK), .Q(net479418), .QN(
        n18112) );
  DFF_X1 \REGISTERS_reg[11][7]  ( .D(n3471), .CK(CLK), .Q(net479417), .QN(
        n18111) );
  DFF_X1 \REGISTERS_reg[11][6]  ( .D(n3470), .CK(CLK), .Q(net479416), .QN(
        n18110) );
  DFF_X1 \REGISTERS_reg[11][5]  ( .D(n3469), .CK(CLK), .Q(net479415), .QN(
        n18109) );
  DFF_X1 \REGISTERS_reg[11][4]  ( .D(n3468), .CK(CLK), .Q(net479414), .QN(
        n18085) );
  DFF_X1 \REGISTERS_reg[11][3]  ( .D(n3467), .CK(CLK), .Q(net479413), .QN(
        n18108) );
  DFF_X1 \REGISTERS_reg[11][2]  ( .D(n3466), .CK(CLK), .Q(net479412), .QN(
        n18084) );
  DFF_X1 \REGISTERS_reg[11][1]  ( .D(n3465), .CK(CLK), .Q(net479411), .QN(
        n18107) );
  DFF_X1 \REGISTERS_reg[11][0]  ( .D(n3464), .CK(CLK), .Q(net479410), .QN(
        n18106) );
  DFF_X1 \REGISTERS_reg[12][31]  ( .D(n3463), .CK(CLK), .Q(net591690), .QN(
        n18007) );
  DFF_X1 \REGISTERS_reg[12][30]  ( .D(n3462), .CK(CLK), .Q(net591689), .QN(
        n18006) );
  DFF_X1 \REGISTERS_reg[12][29]  ( .D(n3461), .CK(CLK), .Q(net591688), .QN(
        n18005) );
  DFF_X1 \REGISTERS_reg[12][28]  ( .D(n3460), .CK(CLK), .Q(net591687), .QN(
        n18004) );
  DFF_X1 \REGISTERS_reg[12][27]  ( .D(n3459), .CK(CLK), .Q(net591686), .QN(
        n18003) );
  DFF_X1 \REGISTERS_reg[12][26]  ( .D(n3458), .CK(CLK), .Q(net591685), .QN(
        n18002) );
  DFF_X1 \REGISTERS_reg[12][25]  ( .D(n3457), .CK(CLK), .Q(net591684), .QN(
        n18001) );
  DFF_X1 \REGISTERS_reg[12][24]  ( .D(n3456), .CK(CLK), .Q(net591683), .QN(
        n18000) );
  DFF_X1 \REGISTERS_reg[12][23]  ( .D(n3455), .CK(CLK), .Q(net591682), .QN(
        n18042) );
  DFF_X1 \REGISTERS_reg[12][22]  ( .D(n3454), .CK(CLK), .Q(net591681), .QN(
        n18041) );
  DFF_X1 \REGISTERS_reg[12][21]  ( .D(n3453), .CK(CLK), .Q(net591680), .QN(
        n18040) );
  DFF_X1 \REGISTERS_reg[12][20]  ( .D(n3452), .CK(CLK), .Q(net591679), .QN(
        n18039) );
  DFF_X1 \REGISTERS_reg[12][19]  ( .D(n3451), .CK(CLK), .Q(net591678), .QN(
        n18038) );
  DFF_X1 \REGISTERS_reg[12][18]  ( .D(n3450), .CK(CLK), .Q(net591677), .QN(
        n18037) );
  DFF_X1 \REGISTERS_reg[12][17]  ( .D(n3449), .CK(CLK), .Q(net591676), .QN(
        n18036) );
  DFF_X1 \REGISTERS_reg[12][16]  ( .D(n3448), .CK(CLK), .Q(net591675), .QN(
        n18035) );
  DFF_X1 \REGISTERS_reg[12][15]  ( .D(n3447), .CK(CLK), .Q(net591674), .QN(
        n18034) );
  DFF_X1 \REGISTERS_reg[12][14]  ( .D(n3446), .CK(CLK), .Q(net591673), .QN(
        n18033) );
  DFF_X1 \REGISTERS_reg[12][13]  ( .D(n3445), .CK(CLK), .Q(net591672), .QN(
        n18032) );
  DFF_X1 \REGISTERS_reg[12][12]  ( .D(n3444), .CK(CLK), .Q(net591671), .QN(
        n18031) );
  DFF_X1 \REGISTERS_reg[12][11]  ( .D(n3443), .CK(CLK), .Q(net591670), .QN(
        n18030) );
  DFF_X1 \REGISTERS_reg[12][10]  ( .D(n3442), .CK(CLK), .Q(net591669), .QN(
        n18029) );
  DFF_X1 \REGISTERS_reg[12][9]  ( .D(n3441), .CK(CLK), .Q(net591668), .QN(
        n18028) );
  DFF_X1 \REGISTERS_reg[12][8]  ( .D(n3440), .CK(CLK), .Q(net591667), .QN(
        n18027) );
  DFF_X1 \REGISTERS_reg[12][7]  ( .D(n3439), .CK(CLK), .Q(net591666), .QN(
        n18026) );
  DFF_X1 \REGISTERS_reg[12][6]  ( .D(n3438), .CK(CLK), .Q(net591665), .QN(
        n18025) );
  DFF_X1 \REGISTERS_reg[12][5]  ( .D(n3437), .CK(CLK), .Q(net591664), .QN(
        n18024) );
  DFF_X1 \REGISTERS_reg[12][4]  ( .D(n3436), .CK(CLK), .Q(net591663), .QN(
        n18018) );
  DFF_X1 \REGISTERS_reg[12][3]  ( .D(n3435), .CK(CLK), .Q(net591662), .QN(
        n18023) );
  DFF_X1 \REGISTERS_reg[12][2]  ( .D(n3434), .CK(CLK), .Q(net591661), .QN(
        n18022) );
  DFF_X1 \REGISTERS_reg[12][1]  ( .D(n3433), .CK(CLK), .Q(net591660), .QN(
        n18017) );
  DFF_X1 \REGISTERS_reg[12][0]  ( .D(n3432), .CK(CLK), .Q(net591659), .QN(
        n18016) );
  DFF_X1 \REGISTERS_reg[13][31]  ( .D(n3431), .CK(CLK), .Q(net479408), .QN(
        n18167) );
  DFF_X1 \REGISTERS_reg[13][30]  ( .D(n3430), .CK(CLK), .Q(net479407), .QN(
        n18166) );
  DFF_X1 \REGISTERS_reg[13][29]  ( .D(n3429), .CK(CLK), .Q(net479406), .QN(
        n18165) );
  DFF_X1 \REGISTERS_reg[13][28]  ( .D(n3428), .CK(CLK), .Q(net479405), .QN(
        n18164) );
  DFF_X1 \REGISTERS_reg[13][27]  ( .D(n3427), .CK(CLK), .Q(net479404), .QN(
        n18163) );
  DFF_X1 \REGISTERS_reg[13][26]  ( .D(n3426), .CK(CLK), .Q(net479403), .QN(
        n18162) );
  DFF_X1 \REGISTERS_reg[13][25]  ( .D(n3425), .CK(CLK), .Q(net479402), .QN(
        n18161) );
  DFF_X1 \REGISTERS_reg[13][24]  ( .D(n3424), .CK(CLK), .Q(net479401), .QN(
        n18160) );
  DFF_X1 \REGISTERS_reg[13][23]  ( .D(n3423), .CK(CLK), .Q(net479400), .QN(
        n18191) );
  DFF_X1 \REGISTERS_reg[13][22]  ( .D(n3422), .CK(CLK), .Q(net479399), .QN(
        n18190) );
  DFF_X1 \REGISTERS_reg[13][21]  ( .D(n3421), .CK(CLK), .Q(net479398), .QN(
        n18189) );
  DFF_X1 \REGISTERS_reg[13][20]  ( .D(n3420), .CK(CLK), .Q(net479397), .QN(
        n18188) );
  DFF_X1 \REGISTERS_reg[13][19]  ( .D(n3419), .CK(CLK), .Q(net479396), .QN(
        n18187) );
  DFF_X1 \REGISTERS_reg[13][18]  ( .D(n3418), .CK(CLK), .Q(net479395), .QN(
        n18186) );
  DFF_X1 \REGISTERS_reg[13][17]  ( .D(n3417), .CK(CLK), .Q(net479394), .QN(
        n18185) );
  DFF_X1 \REGISTERS_reg[13][16]  ( .D(n3416), .CK(CLK), .Q(net479393), .QN(
        n18184) );
  DFF_X1 \REGISTERS_reg[13][15]  ( .D(n3415), .CK(CLK), .Q(net479392), .QN(
        n18183) );
  DFF_X1 \REGISTERS_reg[13][14]  ( .D(n3414), .CK(CLK), .Q(net479391), .QN(
        n18182) );
  DFF_X1 \REGISTERS_reg[13][13]  ( .D(n3413), .CK(CLK), .Q(net479390), .QN(
        n18181) );
  DFF_X1 \REGISTERS_reg[13][12]  ( .D(n3412), .CK(CLK), .Q(net479389), .QN(
        n18180) );
  DFF_X1 \REGISTERS_reg[13][11]  ( .D(n3411), .CK(CLK), .Q(net479388), .QN(
        n18179) );
  DFF_X1 \REGISTERS_reg[13][10]  ( .D(n3410), .CK(CLK), .Q(net479387), .QN(
        n18178) );
  DFF_X1 \REGISTERS_reg[13][9]  ( .D(n3409), .CK(CLK), .Q(net479386), .QN(
        n18177) );
  DFF_X1 \REGISTERS_reg[13][8]  ( .D(n3408), .CK(CLK), .Q(net479385), .QN(
        n18176) );
  DFF_X1 \REGISTERS_reg[13][7]  ( .D(n3407), .CK(CLK), .Q(net479384), .QN(
        n18175) );
  DFF_X1 \REGISTERS_reg[13][6]  ( .D(n3406), .CK(CLK), .Q(net479383), .QN(
        n18174) );
  DFF_X1 \REGISTERS_reg[13][5]  ( .D(n3405), .CK(CLK), .Q(net479382), .QN(
        n18173) );
  DFF_X1 \REGISTERS_reg[13][4]  ( .D(n3404), .CK(CLK), .Q(net479381), .QN(
        n18169) );
  DFF_X1 \REGISTERS_reg[13][3]  ( .D(n3403), .CK(CLK), .Q(net479380), .QN(
        n18172) );
  DFF_X1 \REGISTERS_reg[13][2]  ( .D(n3402), .CK(CLK), .Q(net479379), .QN(
        n18171) );
  DFF_X1 \REGISTERS_reg[13][1]  ( .D(n3401), .CK(CLK), .Q(net479378), .QN(
        n18168) );
  DFF_X1 \REGISTERS_reg[13][0]  ( .D(n3400), .CK(CLK), .Q(net479377), .QN(
        n18170) );
  DFF_X1 \REGISTERS_reg[14][31]  ( .D(n3399), .CK(CLK), .QN(n17847) );
  DFF_X1 \REGISTERS_reg[14][30]  ( .D(n3398), .CK(CLK), .QN(n17846) );
  DFF_X1 \REGISTERS_reg[14][29]  ( .D(n3397), .CK(CLK), .QN(n17845) );
  DFF_X1 \REGISTERS_reg[14][28]  ( .D(n3396), .CK(CLK), .QN(n17844) );
  DFF_X1 \REGISTERS_reg[14][27]  ( .D(n3395), .CK(CLK), .QN(n17843) );
  DFF_X1 \REGISTERS_reg[14][26]  ( .D(n3394), .CK(CLK), .QN(n17842) );
  DFF_X1 \REGISTERS_reg[14][25]  ( .D(n3393), .CK(CLK), .QN(n17841) );
  DFF_X1 \REGISTERS_reg[14][24]  ( .D(n3392), .CK(CLK), .QN(n17840) );
  DFF_X1 \REGISTERS_reg[14][23]  ( .D(n3391), .CK(CLK), .QN(n17871) );
  DFF_X1 \REGISTERS_reg[14][22]  ( .D(n3390), .CK(CLK), .QN(n17870) );
  DFF_X1 \REGISTERS_reg[14][21]  ( .D(n3389), .CK(CLK), .QN(n17869) );
  DFF_X1 \REGISTERS_reg[14][20]  ( .D(n3388), .CK(CLK), .QN(n17868) );
  DFF_X1 \REGISTERS_reg[14][19]  ( .D(n3387), .CK(CLK), .QN(n17867) );
  DFF_X1 \REGISTERS_reg[14][18]  ( .D(n3386), .CK(CLK), .QN(n17866) );
  DFF_X1 \REGISTERS_reg[14][17]  ( .D(n3385), .CK(CLK), .QN(n17865) );
  DFF_X1 \REGISTERS_reg[14][16]  ( .D(n3384), .CK(CLK), .QN(n17864) );
  DFF_X1 \REGISTERS_reg[14][15]  ( .D(n3383), .CK(CLK), .QN(n17863) );
  DFF_X1 \REGISTERS_reg[14][14]  ( .D(n3382), .CK(CLK), .QN(n17862) );
  DFF_X1 \REGISTERS_reg[14][13]  ( .D(n3381), .CK(CLK), .QN(n17861) );
  DFF_X1 \REGISTERS_reg[14][12]  ( .D(n3380), .CK(CLK), .QN(n17860) );
  DFF_X1 \REGISTERS_reg[14][11]  ( .D(n3379), .CK(CLK), .QN(n17859) );
  DFF_X1 \REGISTERS_reg[14][10]  ( .D(n3378), .CK(CLK), .QN(n17858) );
  DFF_X1 \REGISTERS_reg[14][9]  ( .D(n3377), .CK(CLK), .QN(n17857) );
  DFF_X1 \REGISTERS_reg[14][8]  ( .D(n3376), .CK(CLK), .QN(n17856) );
  DFF_X1 \REGISTERS_reg[14][7]  ( .D(n3375), .CK(CLK), .QN(n17855) );
  DFF_X1 \REGISTERS_reg[14][6]  ( .D(n3374), .CK(CLK), .QN(n17854) );
  DFF_X1 \REGISTERS_reg[14][5]  ( .D(n3373), .CK(CLK), .QN(n17853) );
  DFF_X1 \REGISTERS_reg[14][4]  ( .D(n3372), .CK(CLK), .QN(n17852) );
  DFF_X1 \REGISTERS_reg[14][3]  ( .D(n3371), .CK(CLK), .QN(n17851) );
  DFF_X1 \REGISTERS_reg[14][2]  ( .D(n3370), .CK(CLK), .QN(n17850) );
  DFF_X1 \REGISTERS_reg[14][1]  ( .D(n3369), .CK(CLK), .QN(n17849) );
  DFF_X1 \REGISTERS_reg[14][0]  ( .D(n3368), .CK(CLK), .QN(n17848) );
  DFF_X1 \REGISTERS_reg[15][31]  ( .D(n3367), .CK(CLK), .Q(net535499), .QN(
        n18237) );
  DFF_X1 \REGISTERS_reg[15][30]  ( .D(n3366), .CK(CLK), .Q(net535498), .QN(
        n18236) );
  DFF_X1 \REGISTERS_reg[15][29]  ( .D(n3365), .CK(CLK), .Q(net535497), .QN(
        n18235) );
  DFF_X1 \REGISTERS_reg[15][28]  ( .D(n3364), .CK(CLK), .Q(net535496), .QN(
        n18234) );
  DFF_X1 \REGISTERS_reg[15][27]  ( .D(n3363), .CK(CLK), .Q(net535495), .QN(
        n18233) );
  DFF_X1 \REGISTERS_reg[15][26]  ( .D(n3362), .CK(CLK), .Q(net535494), .QN(
        n18232) );
  DFF_X1 \REGISTERS_reg[15][25]  ( .D(n3361), .CK(CLK), .Q(net535493), .QN(
        n18231) );
  DFF_X1 \REGISTERS_reg[15][24]  ( .D(n3360), .CK(CLK), .Q(net535492), .QN(
        n18230) );
  DFF_X1 \REGISTERS_reg[15][23]  ( .D(n3359), .CK(CLK), .Q(net535491), .QN(
        n18253) );
  DFF_X1 \REGISTERS_reg[15][22]  ( .D(n3358), .CK(CLK), .Q(net535490), .QN(
        n18252) );
  DFF_X1 \REGISTERS_reg[15][21]  ( .D(n3357), .CK(CLK), .Q(net535489), .QN(
        n18251) );
  DFF_X1 \REGISTERS_reg[15][20]  ( .D(n3356), .CK(CLK), .Q(net535488), .QN(
        n18250) );
  DFF_X1 \REGISTERS_reg[15][19]  ( .D(n3355), .CK(CLK), .Q(net535487), .QN(
        n18249) );
  DFF_X1 \REGISTERS_reg[15][18]  ( .D(n3354), .CK(CLK), .Q(net535486), .QN(
        n18248) );
  DFF_X1 \REGISTERS_reg[15][17]  ( .D(n3353), .CK(CLK), .Q(net535485), .QN(
        n18247) );
  DFF_X1 \REGISTERS_reg[15][16]  ( .D(n3352), .CK(CLK), .Q(net535484), .QN(
        n18246) );
  DFF_X1 \REGISTERS_reg[15][15]  ( .D(n3351), .CK(CLK), .Q(net535483), .QN(
        n18245) );
  DFF_X1 \REGISTERS_reg[15][14]  ( .D(n3350), .CK(CLK), .Q(net535482), .QN(
        n18244) );
  DFF_X1 \REGISTERS_reg[15][13]  ( .D(n3349), .CK(CLK), .Q(net535481), .QN(
        n18243) );
  DFF_X1 \REGISTERS_reg[15][12]  ( .D(n3348), .CK(CLK), .Q(net535480), .QN(
        n18242) );
  DFF_X1 \REGISTERS_reg[15][11]  ( .D(n3347), .CK(CLK), .Q(net535479), .QN(
        n18241) );
  DFF_X1 \REGISTERS_reg[15][10]  ( .D(n3346), .CK(CLK), .Q(net535478), .QN(
        n18240) );
  DFF_X1 \REGISTERS_reg[15][9]  ( .D(n3345), .CK(CLK), .Q(net535477), .QN(
        n18239) );
  DFF_X1 \REGISTERS_reg[15][8]  ( .D(n3344), .CK(CLK), .Q(net535476), .QN(
        n18238) );
  DFF_X1 \REGISTERS_reg[15][7]  ( .D(n3343), .CK(CLK), .Q(net535475), .QN(
        n18229) );
  DFF_X1 \REGISTERS_reg[15][6]  ( .D(n3342), .CK(CLK), .Q(net535474), .QN(
        n18228) );
  DFF_X1 \REGISTERS_reg[15][5]  ( .D(n3341), .CK(CLK), .Q(net535473), .QN(
        n18227) );
  DFF_X1 \REGISTERS_reg[15][4]  ( .D(n3340), .CK(CLK), .Q(net535472), .QN(
        n18287) );
  DFF_X1 \REGISTERS_reg[15][3]  ( .D(n3339), .CK(CLK), .Q(net535471), .QN(
        n18226) );
  DFF_X1 \REGISTERS_reg[15][2]  ( .D(n3338), .CK(CLK), .Q(net535470), .QN(
        n18225) );
  DFF_X1 \REGISTERS_reg[15][1]  ( .D(n3337), .CK(CLK), .Q(net535469), .QN(
        n18224) );
  DFF_X1 \REGISTERS_reg[15][0]  ( .D(n3336), .CK(CLK), .Q(net535468), .QN(
        n18223) );
  DFF_X1 \REGISTERS_reg[16][31]  ( .D(n3335), .CK(CLK), .Q(net591658), .QN(
        n18071) );
  DFF_X1 \REGISTERS_reg[16][30]  ( .D(n3334), .CK(CLK), .Q(net591657), .QN(
        n18070) );
  DFF_X1 \REGISTERS_reg[16][29]  ( .D(n3333), .CK(CLK), .Q(net591656), .QN(
        n18069) );
  DFF_X1 \REGISTERS_reg[16][28]  ( .D(n3332), .CK(CLK), .Q(net591655), .QN(
        n18068) );
  DFF_X1 \REGISTERS_reg[16][27]  ( .D(n3331), .CK(CLK), .Q(net591654), .QN(
        n18067) );
  DFF_X1 \REGISTERS_reg[16][26]  ( .D(n3330), .CK(CLK), .Q(net591653), .QN(
        n18066) );
  DFF_X1 \REGISTERS_reg[16][25]  ( .D(n3329), .CK(CLK), .Q(net591652), .QN(
        n18065) );
  DFF_X1 \REGISTERS_reg[16][24]  ( .D(n3328), .CK(CLK), .Q(net591651), .QN(
        n18064) );
  DFF_X1 \REGISTERS_reg[16][23]  ( .D(n3327), .CK(CLK), .Q(net591650), .QN(
        n18105) );
  DFF_X1 \REGISTERS_reg[16][22]  ( .D(n3326), .CK(CLK), .Q(net591649), .QN(
        n18104) );
  DFF_X1 \REGISTERS_reg[16][21]  ( .D(n3325), .CK(CLK), .Q(net591648), .QN(
        n18103) );
  DFF_X1 \REGISTERS_reg[16][20]  ( .D(n3324), .CK(CLK), .Q(net591647), .QN(
        n18102) );
  DFF_X1 \REGISTERS_reg[16][19]  ( .D(n3323), .CK(CLK), .Q(net591646), .QN(
        n18101) );
  DFF_X1 \REGISTERS_reg[16][18]  ( .D(n3322), .CK(CLK), .Q(net591645), .QN(
        n18100) );
  DFF_X1 \REGISTERS_reg[16][17]  ( .D(n3321), .CK(CLK), .Q(net591644), .QN(
        n18099) );
  DFF_X1 \REGISTERS_reg[16][16]  ( .D(n3320), .CK(CLK), .Q(net591643), .QN(
        n18098) );
  DFF_X1 \REGISTERS_reg[16][15]  ( .D(n3319), .CK(CLK), .Q(net591642), .QN(
        n18097) );
  DFF_X1 \REGISTERS_reg[16][14]  ( .D(n3318), .CK(CLK), .Q(net591641), .QN(
        n18096) );
  DFF_X1 \REGISTERS_reg[16][13]  ( .D(n3317), .CK(CLK), .Q(net591640), .QN(
        n18095) );
  DFF_X1 \REGISTERS_reg[16][12]  ( .D(n3316), .CK(CLK), .Q(net591639), .QN(
        n18094) );
  DFF_X1 \REGISTERS_reg[16][11]  ( .D(n3315), .CK(CLK), .Q(net591638), .QN(
        n18093) );
  DFF_X1 \REGISTERS_reg[16][10]  ( .D(n3314), .CK(CLK), .Q(net591637), .QN(
        n18092) );
  DFF_X1 \REGISTERS_reg[16][9]  ( .D(n3313), .CK(CLK), .Q(net591636), .QN(
        n18091) );
  DFF_X1 \REGISTERS_reg[16][8]  ( .D(n3312), .CK(CLK), .Q(net591635), .QN(
        n18090) );
  DFF_X1 \REGISTERS_reg[16][7]  ( .D(n3311), .CK(CLK), .Q(net591634), .QN(
        n18089) );
  DFF_X1 \REGISTERS_reg[16][6]  ( .D(n3310), .CK(CLK), .Q(net591633), .QN(
        n18088) );
  DFF_X1 \REGISTERS_reg[16][5]  ( .D(n3309), .CK(CLK), .Q(net591632), .QN(
        n18087) );
  DFF_X1 \REGISTERS_reg[16][4]  ( .D(n3308), .CK(CLK), .Q(net591631), .QN(
        n18086) );
  DFF_X1 \REGISTERS_reg[16][3]  ( .D(n3307), .CK(CLK), .Q(net591630), .QN(
        n18083) );
  DFF_X1 \REGISTERS_reg[16][2]  ( .D(n3306), .CK(CLK), .Q(net591629), .QN(
        n18082) );
  DFF_X1 \REGISTERS_reg[16][1]  ( .D(n3305), .CK(CLK), .Q(net591628), .QN(
        n18081) );
  DFF_X1 \REGISTERS_reg[16][0]  ( .D(n3304), .CK(CLK), .Q(net591627), .QN(
        n18080) );
  DFF_X1 \REGISTERS_reg[17][31]  ( .D(n3303), .CK(CLK), .Q(net423205), .QN(
        n17750) );
  DFF_X1 \REGISTERS_reg[17][30]  ( .D(n3302), .CK(CLK), .Q(net423204), .QN(
        n17749) );
  DFF_X1 \REGISTERS_reg[17][29]  ( .D(n3301), .CK(CLK), .Q(net423203), .QN(
        n17748) );
  DFF_X1 \REGISTERS_reg[17][28]  ( .D(n3300), .CK(CLK), .Q(net423202), .QN(
        n17747) );
  DFF_X1 \REGISTERS_reg[17][27]  ( .D(n3299), .CK(CLK), .Q(net423201), .QN(
        n17746) );
  DFF_X1 \REGISTERS_reg[17][26]  ( .D(n3298), .CK(CLK), .Q(net423200), .QN(
        n17745) );
  DFF_X1 \REGISTERS_reg[17][25]  ( .D(n3297), .CK(CLK), .Q(net423199), .QN(
        n17744) );
  DFF_X1 \REGISTERS_reg[17][24]  ( .D(n3296), .CK(CLK), .Q(net423198), .QN(
        n17743) );
  DFF_X1 \REGISTERS_reg[17][23]  ( .D(n3295), .CK(CLK), .Q(net423197), .QN(
        n17774) );
  DFF_X1 \REGISTERS_reg[17][22]  ( .D(n3294), .CK(CLK), .Q(net423196), .QN(
        n17773) );
  DFF_X1 \REGISTERS_reg[17][21]  ( .D(n3293), .CK(CLK), .Q(net423195), .QN(
        n17772) );
  DFF_X1 \REGISTERS_reg[17][20]  ( .D(n3292), .CK(CLK), .Q(net423194), .QN(
        n17771) );
  DFF_X1 \REGISTERS_reg[17][19]  ( .D(n3291), .CK(CLK), .Q(net423193), .QN(
        n17770) );
  DFF_X1 \REGISTERS_reg[17][18]  ( .D(n3290), .CK(CLK), .Q(net423192), .QN(
        n17769) );
  DFF_X1 \REGISTERS_reg[17][17]  ( .D(n3289), .CK(CLK), .Q(net423191), .QN(
        n17768) );
  DFF_X1 \REGISTERS_reg[17][16]  ( .D(n3288), .CK(CLK), .Q(net423190), .QN(
        n17767) );
  DFF_X1 \REGISTERS_reg[17][15]  ( .D(n3287), .CK(CLK), .Q(net423189), .QN(
        n17766) );
  DFF_X1 \REGISTERS_reg[17][14]  ( .D(n3286), .CK(CLK), .Q(net423188), .QN(
        n17765) );
  DFF_X1 \REGISTERS_reg[17][13]  ( .D(n3285), .CK(CLK), .Q(net423187), .QN(
        n17764) );
  DFF_X1 \REGISTERS_reg[17][12]  ( .D(n3284), .CK(CLK), .Q(net423186), .QN(
        n17763) );
  DFF_X1 \REGISTERS_reg[17][11]  ( .D(n3283), .CK(CLK), .Q(net423185), .QN(
        n17762) );
  DFF_X1 \REGISTERS_reg[17][10]  ( .D(n3282), .CK(CLK), .Q(net423184), .QN(
        n17761) );
  DFF_X1 \REGISTERS_reg[17][9]  ( .D(n3281), .CK(CLK), .Q(net423183), .QN(
        n17760) );
  DFF_X1 \REGISTERS_reg[17][8]  ( .D(n3280), .CK(CLK), .Q(net423182), .QN(
        n17759) );
  DFF_X1 \REGISTERS_reg[17][7]  ( .D(n3279), .CK(CLK), .Q(net423181), .QN(
        n17758) );
  DFF_X1 \REGISTERS_reg[17][6]  ( .D(n3278), .CK(CLK), .Q(net423180), .QN(
        n17757) );
  DFF_X1 \REGISTERS_reg[17][5]  ( .D(n3277), .CK(CLK), .Q(net423179), .QN(
        n17756) );
  DFF_X1 \REGISTERS_reg[17][4]  ( .D(n3276), .CK(CLK), .Q(net423178), .QN(
        n17755) );
  DFF_X1 \REGISTERS_reg[17][3]  ( .D(n3275), .CK(CLK), .Q(net423177), .QN(
        n17753) );
  DFF_X1 \REGISTERS_reg[17][2]  ( .D(n3274), .CK(CLK), .Q(net423176), .QN(
        n17752) );
  DFF_X1 \REGISTERS_reg[17][1]  ( .D(n3273), .CK(CLK), .Q(net423175), .QN(
        n17751) );
  DFF_X1 \REGISTERS_reg[17][0]  ( .D(n3272), .CK(CLK), .Q(net423174), .QN(
        n17754) );
  DFF_X1 \REGISTERS_reg[18][31]  ( .D(n3271), .CK(CLK), .Q(net367046), .QN(
        n17879) );
  DFF_X1 \REGISTERS_reg[18][30]  ( .D(n3270), .CK(CLK), .Q(net367045), .QN(
        n17878) );
  DFF_X1 \REGISTERS_reg[18][29]  ( .D(n3269), .CK(CLK), .Q(net367044), .QN(
        n17877) );
  DFF_X1 \REGISTERS_reg[18][28]  ( .D(n3268), .CK(CLK), .Q(net367043), .QN(
        n17876) );
  DFF_X1 \REGISTERS_reg[18][27]  ( .D(n3267), .CK(CLK), .Q(net367042), .QN(
        n17875) );
  DFF_X1 \REGISTERS_reg[18][26]  ( .D(n3266), .CK(CLK), .Q(net367041), .QN(
        n17874) );
  DFF_X1 \REGISTERS_reg[18][25]  ( .D(n3265), .CK(CLK), .Q(net367040), .QN(
        n17873) );
  DFF_X1 \REGISTERS_reg[18][24]  ( .D(n3264), .CK(CLK), .Q(net367039), .QN(
        n17872) );
  DFF_X1 \REGISTERS_reg[18][23]  ( .D(n3263), .CK(CLK), .Q(net367038), .QN(
        n17903) );
  DFF_X1 \REGISTERS_reg[18][22]  ( .D(n3262), .CK(CLK), .Q(net367037), .QN(
        n17902) );
  DFF_X1 \REGISTERS_reg[18][21]  ( .D(n3261), .CK(CLK), .Q(net367036), .QN(
        n17901) );
  DFF_X1 \REGISTERS_reg[18][20]  ( .D(n3260), .CK(CLK), .Q(net367035), .QN(
        n17900) );
  DFF_X1 \REGISTERS_reg[18][19]  ( .D(n3259), .CK(CLK), .Q(net367034), .QN(
        n17899) );
  DFF_X1 \REGISTERS_reg[18][18]  ( .D(n3258), .CK(CLK), .Q(net367033), .QN(
        n17898) );
  DFF_X1 \REGISTERS_reg[18][17]  ( .D(n3257), .CK(CLK), .Q(net367032), .QN(
        n17897) );
  DFF_X1 \REGISTERS_reg[18][16]  ( .D(n3256), .CK(CLK), .Q(net367031), .QN(
        n17896) );
  DFF_X1 \REGISTERS_reg[18][15]  ( .D(n3255), .CK(CLK), .Q(net367030), .QN(
        n17895) );
  DFF_X1 \REGISTERS_reg[18][14]  ( .D(n3254), .CK(CLK), .Q(net367029), .QN(
        n17894) );
  DFF_X1 \REGISTERS_reg[18][13]  ( .D(n3253), .CK(CLK), .Q(net367028), .QN(
        n17893) );
  DFF_X1 \REGISTERS_reg[18][12]  ( .D(n3252), .CK(CLK), .Q(net367027), .QN(
        n17892) );
  DFF_X1 \REGISTERS_reg[18][11]  ( .D(n3251), .CK(CLK), .Q(net367026), .QN(
        n17891) );
  DFF_X1 \REGISTERS_reg[18][10]  ( .D(n3250), .CK(CLK), .Q(net367025), .QN(
        n17890) );
  DFF_X1 \REGISTERS_reg[18][9]  ( .D(n3249), .CK(CLK), .Q(net367024), .QN(
        n17889) );
  DFF_X1 \REGISTERS_reg[18][8]  ( .D(n3248), .CK(CLK), .Q(net367023), .QN(
        n17888) );
  DFF_X1 \REGISTERS_reg[18][7]  ( .D(n3247), .CK(CLK), .Q(net367022), .QN(
        n17887) );
  DFF_X1 \REGISTERS_reg[18][6]  ( .D(n3246), .CK(CLK), .Q(net367021), .QN(
        n17886) );
  DFF_X1 \REGISTERS_reg[18][5]  ( .D(n3245), .CK(CLK), .Q(net367020), .QN(
        n17885) );
  DFF_X1 \REGISTERS_reg[18][4]  ( .D(n3244), .CK(CLK), .Q(net367019), .QN(
        n17884) );
  DFF_X1 \REGISTERS_reg[18][3]  ( .D(n3243), .CK(CLK), .Q(net367018), .QN(
        n17882) );
  DFF_X1 \REGISTERS_reg[18][2]  ( .D(n3242), .CK(CLK), .Q(net367017), .QN(
        n17881) );
  DFF_X1 \REGISTERS_reg[18][1]  ( .D(n3241), .CK(CLK), .Q(net367016), .QN(
        n17883) );
  DFF_X1 \REGISTERS_reg[18][0]  ( .D(n3240), .CK(CLK), .Q(net367015), .QN(
        n17880) );
  DFF_X1 \REGISTERS_reg[19][31]  ( .D(n3239), .CK(CLK), .Q(net479376), .QN(
        n18135) );
  DFF_X1 \REGISTERS_reg[19][30]  ( .D(n3238), .CK(CLK), .Q(net479375), .QN(
        n18134) );
  DFF_X1 \REGISTERS_reg[19][29]  ( .D(n3237), .CK(CLK), .Q(net479374), .QN(
        n18133) );
  DFF_X1 \REGISTERS_reg[19][28]  ( .D(n3236), .CK(CLK), .Q(net479373), .QN(
        n18132) );
  DFF_X1 \REGISTERS_reg[19][27]  ( .D(n3235), .CK(CLK), .Q(net479372), .QN(
        n18131) );
  DFF_X1 \REGISTERS_reg[19][26]  ( .D(n3234), .CK(CLK), .Q(net479371), .QN(
        n18130) );
  DFF_X1 \REGISTERS_reg[19][25]  ( .D(n3233), .CK(CLK), .Q(net479370), .QN(
        n18129) );
  DFF_X1 \REGISTERS_reg[19][24]  ( .D(n3232), .CK(CLK), .Q(net479369), .QN(
        n18128) );
  DFF_X1 \REGISTERS_reg[19][23]  ( .D(n3231), .CK(CLK), .Q(net479368), .QN(
        n18159) );
  DFF_X1 \REGISTERS_reg[19][22]  ( .D(n3230), .CK(CLK), .Q(net479367), .QN(
        n18158) );
  DFF_X1 \REGISTERS_reg[19][21]  ( .D(n3229), .CK(CLK), .Q(net479366), .QN(
        n18157) );
  DFF_X1 \REGISTERS_reg[19][20]  ( .D(n3228), .CK(CLK), .Q(net479365), .QN(
        n18156) );
  DFF_X1 \REGISTERS_reg[19][19]  ( .D(n3227), .CK(CLK), .Q(net479364), .QN(
        n18155) );
  DFF_X1 \REGISTERS_reg[19][18]  ( .D(n3226), .CK(CLK), .Q(net479363), .QN(
        n18154) );
  DFF_X1 \REGISTERS_reg[19][17]  ( .D(n3225), .CK(CLK), .Q(net479362), .QN(
        n18153) );
  DFF_X1 \REGISTERS_reg[19][16]  ( .D(n3224), .CK(CLK), .Q(net479361), .QN(
        n18152) );
  DFF_X1 \REGISTERS_reg[19][15]  ( .D(n3223), .CK(CLK), .Q(net479360), .QN(
        n18151) );
  DFF_X1 \REGISTERS_reg[19][14]  ( .D(n3222), .CK(CLK), .Q(net479359), .QN(
        n18150) );
  DFF_X1 \REGISTERS_reg[19][13]  ( .D(n3221), .CK(CLK), .Q(net479358), .QN(
        n18149) );
  DFF_X1 \REGISTERS_reg[19][12]  ( .D(n3220), .CK(CLK), .Q(net479357), .QN(
        n18148) );
  DFF_X1 \REGISTERS_reg[19][11]  ( .D(n3219), .CK(CLK), .Q(net479356), .QN(
        n18147) );
  DFF_X1 \REGISTERS_reg[19][10]  ( .D(n3218), .CK(CLK), .Q(net479355), .QN(
        n18146) );
  DFF_X1 \REGISTERS_reg[19][9]  ( .D(n3217), .CK(CLK), .Q(net479354), .QN(
        n18145) );
  DFF_X1 \REGISTERS_reg[19][8]  ( .D(n3216), .CK(CLK), .Q(net479353), .QN(
        n18144) );
  DFF_X1 \REGISTERS_reg[19][7]  ( .D(n3215), .CK(CLK), .Q(net479352), .QN(
        n18143) );
  DFF_X1 \REGISTERS_reg[19][6]  ( .D(n3214), .CK(CLK), .Q(net479351), .QN(
        n18142) );
  DFF_X1 \REGISTERS_reg[19][5]  ( .D(n3213), .CK(CLK), .Q(net479350), .QN(
        n18141) );
  DFF_X1 \REGISTERS_reg[19][4]  ( .D(n3212), .CK(CLK), .Q(net479349), .QN(
        n18140) );
  DFF_X1 \REGISTERS_reg[19][3]  ( .D(n3211), .CK(CLK), .Q(net479348), .QN(
        n18137) );
  DFF_X1 \REGISTERS_reg[19][2]  ( .D(n3210), .CK(CLK), .Q(net479347), .QN(
        n18136) );
  DFF_X1 \REGISTERS_reg[19][1]  ( .D(n3209), .CK(CLK), .Q(net479346), .QN(
        n18139) );
  DFF_X1 \REGISTERS_reg[19][0]  ( .D(n3208), .CK(CLK), .Q(net479345), .QN(
        n18138) );
  DFF_X1 \REGISTERS_reg[20][31]  ( .D(n3207), .CK(CLK), .Q(net366982), .QN(
        n18295) );
  DFF_X1 \REGISTERS_reg[20][30]  ( .D(n3206), .CK(CLK), .Q(net366981), .QN(
        n18294) );
  DFF_X1 \REGISTERS_reg[20][29]  ( .D(n3205), .CK(CLK), .Q(net366980), .QN(
        n18293) );
  DFF_X1 \REGISTERS_reg[20][28]  ( .D(n3204), .CK(CLK), .Q(net366979), .QN(
        n18292) );
  DFF_X1 \REGISTERS_reg[20][27]  ( .D(n3203), .CK(CLK), .Q(net366978), .QN(
        n18291) );
  DFF_X1 \REGISTERS_reg[20][26]  ( .D(n3202), .CK(CLK), .Q(net366977), .QN(
        n18290) );
  DFF_X1 \REGISTERS_reg[20][25]  ( .D(n3201), .CK(CLK), .Q(net366976), .QN(
        n18289) );
  DFF_X1 \REGISTERS_reg[20][24]  ( .D(n3200), .CK(CLK), .Q(net366975), .QN(
        n18288) );
  DFF_X1 \REGISTERS_reg[20][23]  ( .D(n3199), .CK(CLK), .Q(net366974), .QN(
        n18319) );
  DFF_X1 \REGISTERS_reg[20][22]  ( .D(n3198), .CK(CLK), .Q(net366973), .QN(
        n18318) );
  DFF_X1 \REGISTERS_reg[20][21]  ( .D(n3197), .CK(CLK), .Q(net366972), .QN(
        n18317) );
  DFF_X1 \REGISTERS_reg[20][20]  ( .D(n3196), .CK(CLK), .Q(net366971), .QN(
        n18316) );
  DFF_X1 \REGISTERS_reg[20][19]  ( .D(n3195), .CK(CLK), .Q(net366970), .QN(
        n18315) );
  DFF_X1 \REGISTERS_reg[20][18]  ( .D(n3194), .CK(CLK), .Q(net366969), .QN(
        n18314) );
  DFF_X1 \REGISTERS_reg[20][17]  ( .D(n3193), .CK(CLK), .Q(net366968), .QN(
        n18313) );
  DFF_X1 \REGISTERS_reg[20][16]  ( .D(n3192), .CK(CLK), .Q(net366967), .QN(
        n18312) );
  DFF_X1 \REGISTERS_reg[20][15]  ( .D(n3191), .CK(CLK), .Q(net366966), .QN(
        n18311) );
  DFF_X1 \REGISTERS_reg[20][14]  ( .D(n3190), .CK(CLK), .Q(net366965), .QN(
        n18310) );
  DFF_X1 \REGISTERS_reg[20][13]  ( .D(n3189), .CK(CLK), .Q(net366964), .QN(
        n18309) );
  DFF_X1 \REGISTERS_reg[20][12]  ( .D(n3188), .CK(CLK), .Q(net366963), .QN(
        n18308) );
  DFF_X1 \REGISTERS_reg[20][11]  ( .D(n3187), .CK(CLK), .Q(net366962), .QN(
        n18307) );
  DFF_X1 \REGISTERS_reg[20][10]  ( .D(n3186), .CK(CLK), .Q(net366961), .QN(
        n18306) );
  DFF_X1 \REGISTERS_reg[20][9]  ( .D(n3185), .CK(CLK), .Q(net366960), .QN(
        n18305) );
  DFF_X1 \REGISTERS_reg[20][8]  ( .D(n3184), .CK(CLK), .Q(net366959), .QN(
        n18304) );
  DFF_X1 \REGISTERS_reg[20][7]  ( .D(n3183), .CK(CLK), .Q(net366958), .QN(
        n18303) );
  DFF_X1 \REGISTERS_reg[20][6]  ( .D(n3182), .CK(CLK), .Q(net366957), .QN(
        n18302) );
  DFF_X1 \REGISTERS_reg[20][5]  ( .D(n3181), .CK(CLK), .Q(net366956), .QN(
        n18301) );
  DFF_X1 \REGISTERS_reg[20][4]  ( .D(n3180), .CK(CLK), .Q(net366955), .QN(
        n18300) );
  DFF_X1 \REGISTERS_reg[20][3]  ( .D(n3179), .CK(CLK), .Q(net366954), .QN(
        n18298) );
  DFF_X1 \REGISTERS_reg[20][2]  ( .D(n3178), .CK(CLK), .Q(net366953), .QN(
        n18299) );
  DFF_X1 \REGISTERS_reg[20][1]  ( .D(n3177), .CK(CLK), .Q(net366952), .QN(
        n18297) );
  DFF_X1 \REGISTERS_reg[20][0]  ( .D(n3176), .CK(CLK), .Q(net366951), .QN(
        n18296) );
  DFF_X1 \REGISTERS_reg[21][31]  ( .D(n3175), .CK(CLK), .QN(n17621) );
  DFF_X1 \REGISTERS_reg[21][30]  ( .D(n3174), .CK(CLK), .QN(n17620) );
  DFF_X1 \REGISTERS_reg[21][29]  ( .D(n3173), .CK(CLK), .QN(n17619) );
  DFF_X1 \REGISTERS_reg[21][28]  ( .D(n3172), .CK(CLK), .QN(n17618) );
  DFF_X1 \REGISTERS_reg[21][27]  ( .D(n3171), .CK(CLK), .QN(n17617) );
  DFF_X1 \REGISTERS_reg[21][26]  ( .D(n3170), .CK(CLK), .QN(n17616) );
  DFF_X1 \REGISTERS_reg[21][25]  ( .D(n3169), .CK(CLK), .QN(n17615) );
  DFF_X1 \REGISTERS_reg[21][24]  ( .D(n3168), .CK(CLK), .QN(n17614) );
  DFF_X1 \REGISTERS_reg[21][23]  ( .D(n3167), .CK(CLK), .QN(n17637) );
  DFF_X1 \REGISTERS_reg[21][22]  ( .D(n3166), .CK(CLK), .QN(n17636) );
  DFF_X1 \REGISTERS_reg[21][21]  ( .D(n3165), .CK(CLK), .QN(n17635) );
  DFF_X1 \REGISTERS_reg[21][20]  ( .D(n3164), .CK(CLK), .QN(n17634) );
  DFF_X1 \REGISTERS_reg[21][19]  ( .D(n3163), .CK(CLK), .QN(n17633) );
  DFF_X1 \REGISTERS_reg[21][18]  ( .D(n3162), .CK(CLK), .QN(n17632) );
  DFF_X1 \REGISTERS_reg[21][17]  ( .D(n3161), .CK(CLK), .QN(n17631) );
  DFF_X1 \REGISTERS_reg[21][16]  ( .D(n3160), .CK(CLK), .QN(n17630) );
  DFF_X1 \REGISTERS_reg[21][15]  ( .D(n3159), .CK(CLK), .QN(n17629) );
  DFF_X1 \REGISTERS_reg[21][14]  ( .D(n3158), .CK(CLK), .QN(n17628) );
  DFF_X1 \REGISTERS_reg[21][13]  ( .D(n3157), .CK(CLK), .QN(n17627) );
  DFF_X1 \REGISTERS_reg[21][12]  ( .D(n3156), .CK(CLK), .QN(n17626) );
  DFF_X1 \REGISTERS_reg[21][11]  ( .D(n3155), .CK(CLK), .QN(n17625) );
  DFF_X1 \REGISTERS_reg[21][10]  ( .D(n3154), .CK(CLK), .QN(n17624) );
  DFF_X1 \REGISTERS_reg[21][9]  ( .D(n3153), .CK(CLK), .QN(n17623) );
  DFF_X1 \REGISTERS_reg[21][8]  ( .D(n3152), .CK(CLK), .QN(n17622) );
  DFF_X1 \REGISTERS_reg[21][7]  ( .D(n3151), .CK(CLK), .QN(n17676) );
  DFF_X1 \REGISTERS_reg[21][6]  ( .D(n3150), .CK(CLK), .QN(n17675) );
  DFF_X1 \REGISTERS_reg[21][5]  ( .D(n3149), .CK(CLK), .QN(n17674) );
  DFF_X1 \REGISTERS_reg[21][4]  ( .D(n3148), .CK(CLK), .QN(n17673) );
  DFF_X1 \REGISTERS_reg[21][3]  ( .D(n3147), .CK(CLK), .QN(n17672) );
  DFF_X1 \REGISTERS_reg[21][2]  ( .D(n3146), .CK(CLK), .QN(n17671) );
  DFF_X1 \REGISTERS_reg[21][1]  ( .D(n3145), .CK(CLK), .QN(n17670) );
  DFF_X1 \REGISTERS_reg[21][0]  ( .D(n3144), .CK(CLK), .QN(n17669) );
  DFF_X1 \REGISTERS_reg[22][31]  ( .D(n3143), .CK(CLK), .Q(net535467), .QN(
        n17782) );
  DFF_X1 \REGISTERS_reg[22][30]  ( .D(n3142), .CK(CLK), .Q(net535466), .QN(
        n17781) );
  DFF_X1 \REGISTERS_reg[22][29]  ( .D(n3141), .CK(CLK), .Q(net535465), .QN(
        n17780) );
  DFF_X1 \REGISTERS_reg[22][28]  ( .D(n3140), .CK(CLK), .Q(net535464), .QN(
        n17779) );
  DFF_X1 \REGISTERS_reg[22][27]  ( .D(n3139), .CK(CLK), .Q(net535463), .QN(
        n17778) );
  DFF_X1 \REGISTERS_reg[22][26]  ( .D(n3138), .CK(CLK), .Q(net535462), .QN(
        n17777) );
  DFF_X1 \REGISTERS_reg[22][25]  ( .D(n3137), .CK(CLK), .Q(net535461), .QN(
        n17776) );
  DFF_X1 \REGISTERS_reg[22][24]  ( .D(n3136), .CK(CLK), .Q(net535460), .QN(
        n17775) );
  DFF_X1 \REGISTERS_reg[22][23]  ( .D(n3135), .CK(CLK), .Q(net535459), .QN(
        n17806) );
  DFF_X1 \REGISTERS_reg[22][22]  ( .D(n3134), .CK(CLK), .Q(net535458), .QN(
        n17805) );
  DFF_X1 \REGISTERS_reg[22][21]  ( .D(n3133), .CK(CLK), .Q(net535457), .QN(
        n17804) );
  DFF_X1 \REGISTERS_reg[22][20]  ( .D(n3132), .CK(CLK), .Q(net535456), .QN(
        n17803) );
  DFF_X1 \REGISTERS_reg[22][19]  ( .D(n3131), .CK(CLK), .Q(net535455), .QN(
        n17802) );
  DFF_X1 \REGISTERS_reg[22][18]  ( .D(n3130), .CK(CLK), .Q(net535454), .QN(
        n17801) );
  DFF_X1 \REGISTERS_reg[22][17]  ( .D(n3129), .CK(CLK), .Q(net535453), .QN(
        n17800) );
  DFF_X1 \REGISTERS_reg[22][16]  ( .D(n3128), .CK(CLK), .Q(net535452), .QN(
        n17799) );
  DFF_X1 \REGISTERS_reg[22][15]  ( .D(n3127), .CK(CLK), .Q(net535451), .QN(
        n17798) );
  DFF_X1 \REGISTERS_reg[22][14]  ( .D(n3126), .CK(CLK), .Q(net535450), .QN(
        n17797) );
  DFF_X1 \REGISTERS_reg[22][13]  ( .D(n3125), .CK(CLK), .Q(net535449), .QN(
        n17796) );
  DFF_X1 \REGISTERS_reg[22][12]  ( .D(n3124), .CK(CLK), .Q(net535448), .QN(
        n17795) );
  DFF_X1 \REGISTERS_reg[22][11]  ( .D(n3123), .CK(CLK), .Q(net535447), .QN(
        n17794) );
  DFF_X1 \REGISTERS_reg[22][10]  ( .D(n3122), .CK(CLK), .Q(net535446), .QN(
        n17793) );
  DFF_X1 \REGISTERS_reg[22][9]  ( .D(n3121), .CK(CLK), .Q(net535445), .QN(
        n17792) );
  DFF_X1 \REGISTERS_reg[22][8]  ( .D(n3120), .CK(CLK), .Q(net535444), .QN(
        n17791) );
  DFF_X1 \REGISTERS_reg[22][7]  ( .D(n3119), .CK(CLK), .Q(net535443), .QN(
        n17790) );
  DFF_X1 \REGISTERS_reg[22][6]  ( .D(n3118), .CK(CLK), .Q(net535442), .QN(
        n17789) );
  DFF_X1 \REGISTERS_reg[22][5]  ( .D(n3117), .CK(CLK), .Q(net535441), .QN(
        n17788) );
  DFF_X1 \REGISTERS_reg[22][4]  ( .D(n3116), .CK(CLK), .Q(net535440), .QN(
        n17787) );
  DFF_X1 \REGISTERS_reg[22][3]  ( .D(n3115), .CK(CLK), .Q(net535439), .QN(
        n17784) );
  DFF_X1 \REGISTERS_reg[22][2]  ( .D(n3114), .CK(CLK), .Q(net535438), .QN(
        n17786) );
  DFF_X1 \REGISTERS_reg[22][1]  ( .D(n3113), .CK(CLK), .Q(net535437), .QN(
        n17785) );
  DFF_X1 \REGISTERS_reg[22][0]  ( .D(n3112), .CK(CLK), .Q(net535436), .QN(
        n17783) );
  DFF_X1 \REGISTERS_reg[23][31]  ( .D(n3111), .CK(CLK), .Q(net310533), .QN(
        n18222) );
  DFF_X1 \REGISTERS_reg[23][30]  ( .D(n3110), .CK(CLK), .Q(net310532), .QN(
        n18221) );
  DFF_X1 \REGISTERS_reg[23][29]  ( .D(n3109), .CK(CLK), .Q(net310531), .QN(
        n18220) );
  DFF_X1 \REGISTERS_reg[23][28]  ( .D(n3108), .CK(CLK), .Q(net310530), .QN(
        n18219) );
  DFF_X1 \REGISTERS_reg[23][27]  ( .D(n3107), .CK(CLK), .Q(net310529), .QN(
        n18218) );
  DFF_X1 \REGISTERS_reg[23][26]  ( .D(n3106), .CK(CLK), .Q(net310528), .QN(
        n18217) );
  DFF_X1 \REGISTERS_reg[23][25]  ( .D(n3105), .CK(CLK), .Q(net310527), .QN(
        n18216) );
  DFF_X1 \REGISTERS_reg[23][24]  ( .D(n3104), .CK(CLK), .Q(net310526), .QN(
        n18215) );
  DFF_X1 \REGISTERS_reg[23][23]  ( .D(n3103), .CK(CLK), .Q(net310525), .QN(
        n18214) );
  DFF_X1 \REGISTERS_reg[23][22]  ( .D(n3102), .CK(CLK), .Q(net310524), .QN(
        n18213) );
  DFF_X1 \REGISTERS_reg[23][21]  ( .D(n3101), .CK(CLK), .Q(net310523), .QN(
        n18212) );
  DFF_X1 \REGISTERS_reg[23][20]  ( .D(n3100), .CK(CLK), .Q(net310522), .QN(
        n18211) );
  DFF_X1 \REGISTERS_reg[23][19]  ( .D(n3099), .CK(CLK), .Q(net310521), .QN(
        n18210) );
  DFF_X1 \REGISTERS_reg[23][18]  ( .D(n3098), .CK(CLK), .Q(net310520), .QN(
        n18209) );
  DFF_X1 \REGISTERS_reg[23][17]  ( .D(n3097), .CK(CLK), .Q(net310519), .QN(
        n18208) );
  DFF_X1 \REGISTERS_reg[23][16]  ( .D(n3096), .CK(CLK), .Q(net310518), .QN(
        n18207) );
  DFF_X1 \REGISTERS_reg[23][15]  ( .D(n3095), .CK(CLK), .Q(net310517), .QN(
        n18206) );
  DFF_X1 \REGISTERS_reg[23][14]  ( .D(n3094), .CK(CLK), .Q(net310516), .QN(
        n18205) );
  DFF_X1 \REGISTERS_reg[23][13]  ( .D(n3093), .CK(CLK), .Q(net310515), .QN(
        n18204) );
  DFF_X1 \REGISTERS_reg[23][12]  ( .D(n3092), .CK(CLK), .Q(net310514), .QN(
        n18203) );
  DFF_X1 \REGISTERS_reg[23][11]  ( .D(n3091), .CK(CLK), .Q(net310513), .QN(
        n18202) );
  DFF_X1 \REGISTERS_reg[23][10]  ( .D(n3090), .CK(CLK), .Q(net310512), .QN(
        n18201) );
  DFF_X1 \REGISTERS_reg[23][9]  ( .D(n3089), .CK(CLK), .Q(net310511), .QN(
        n18200) );
  DFF_X1 \REGISTERS_reg[23][8]  ( .D(n3088), .CK(CLK), .Q(net310510), .QN(
        n18199) );
  DFF_X1 \REGISTERS_reg[23][7]  ( .D(n3087), .CK(CLK), .Q(net310509), .QN(
        n18198) );
  DFF_X1 \REGISTERS_reg[23][6]  ( .D(n3086), .CK(CLK), .Q(net310508), .QN(
        n18197) );
  DFF_X1 \REGISTERS_reg[23][5]  ( .D(n3085), .CK(CLK), .Q(net310507), .QN(
        n18196) );
  DFF_X1 \REGISTERS_reg[23][4]  ( .D(n3084), .CK(CLK), .Q(net310506), .QN(
        n18195) );
  DFF_X1 \REGISTERS_reg[23][3]  ( .D(n3083), .CK(CLK), .Q(net310505), .QN(
        n18286) );
  DFF_X1 \REGISTERS_reg[23][2]  ( .D(n3082), .CK(CLK), .Q(net310504), .QN(
        n18194) );
  DFF_X1 \REGISTERS_reg[23][1]  ( .D(n3081), .CK(CLK), .Q(net310503), .QN(
        n18193) );
  DFF_X1 \REGISTERS_reg[23][0]  ( .D(n3080), .CK(CLK), .Q(net310502), .QN(
        n18192) );
  DFF_X1 \REGISTERS_reg[24][31]  ( .D(n3079), .CK(CLK), .QN(n17366) );
  DFF_X1 \REGISTERS_reg[24][30]  ( .D(n3078), .CK(CLK), .QN(n17365) );
  DFF_X1 \REGISTERS_reg[24][29]  ( .D(n3077), .CK(CLK), .QN(n17364) );
  DFF_X1 \REGISTERS_reg[24][28]  ( .D(n3076), .CK(CLK), .QN(n17363) );
  DFF_X1 \REGISTERS_reg[24][27]  ( .D(n3075), .CK(CLK), .QN(n17362) );
  DFF_X1 \REGISTERS_reg[24][26]  ( .D(n3074), .CK(CLK), .QN(n17361) );
  DFF_X1 \REGISTERS_reg[24][25]  ( .D(n3073), .CK(CLK), .QN(n17360) );
  DFF_X1 \REGISTERS_reg[24][24]  ( .D(n3072), .CK(CLK), .QN(n17359) );
  DFF_X1 \REGISTERS_reg[24][23]  ( .D(n3071), .CK(CLK), .QN(n17382) );
  DFF_X1 \REGISTERS_reg[24][22]  ( .D(n3070), .CK(CLK), .QN(n17381) );
  DFF_X1 \REGISTERS_reg[24][21]  ( .D(n3069), .CK(CLK), .QN(n17380) );
  DFF_X1 \REGISTERS_reg[24][20]  ( .D(n3068), .CK(CLK), .QN(n17379) );
  DFF_X1 \REGISTERS_reg[24][19]  ( .D(n3067), .CK(CLK), .QN(n17378) );
  DFF_X1 \REGISTERS_reg[24][18]  ( .D(n3066), .CK(CLK), .QN(n17377) );
  DFF_X1 \REGISTERS_reg[24][17]  ( .D(n3065), .CK(CLK), .QN(n17376) );
  DFF_X1 \REGISTERS_reg[24][16]  ( .D(n3064), .CK(CLK), .QN(n17375) );
  DFF_X1 \REGISTERS_reg[24][15]  ( .D(n3063), .CK(CLK), .QN(n17374) );
  DFF_X1 \REGISTERS_reg[24][14]  ( .D(n3062), .CK(CLK), .QN(n17373) );
  DFF_X1 \REGISTERS_reg[24][13]  ( .D(n3061), .CK(CLK), .QN(n17372) );
  DFF_X1 \REGISTERS_reg[24][12]  ( .D(n3060), .CK(CLK), .QN(n17371) );
  DFF_X1 \REGISTERS_reg[24][11]  ( .D(n3059), .CK(CLK), .QN(n17370) );
  DFF_X1 \REGISTERS_reg[24][10]  ( .D(n3058), .CK(CLK), .QN(n17369) );
  DFF_X1 \REGISTERS_reg[24][9]  ( .D(n3057), .CK(CLK), .QN(n17368) );
  DFF_X1 \REGISTERS_reg[24][8]  ( .D(n3056), .CK(CLK), .QN(n17367) );
  DFF_X1 \REGISTERS_reg[24][7]  ( .D(n3055), .CK(CLK), .QN(n17390) );
  DFF_X1 \REGISTERS_reg[24][6]  ( .D(n3054), .CK(CLK), .QN(n17389) );
  DFF_X1 \REGISTERS_reg[24][5]  ( .D(n3053), .CK(CLK), .QN(n17388) );
  DFF_X1 \REGISTERS_reg[24][4]  ( .D(n3052), .CK(CLK), .QN(n17387) );
  DFF_X1 \REGISTERS_reg[24][3]  ( .D(n3051), .CK(CLK), .QN(n17386) );
  DFF_X1 \REGISTERS_reg[24][2]  ( .D(n3050), .CK(CLK), .QN(n17385) );
  DFF_X1 \REGISTERS_reg[24][1]  ( .D(n3049), .CK(CLK), .QN(n17384) );
  DFF_X1 \REGISTERS_reg[24][0]  ( .D(n3048), .CK(CLK), .QN(n17383) );
  DFF_X1 \REGISTERS_reg[25][31]  ( .D(n3047), .CK(CLK), .Q(net479344), .QN(
        n17911) );
  DFF_X1 \REGISTERS_reg[25][30]  ( .D(n3046), .CK(CLK), .Q(net310500), .QN(
        n17910) );
  DFF_X1 \REGISTERS_reg[25][29]  ( .D(n3045), .CK(CLK), .Q(net310499), .QN(
        n17909) );
  DFF_X1 \REGISTERS_reg[25][28]  ( .D(n3044), .CK(CLK), .Q(net310498), .QN(
        n17908) );
  DFF_X1 \REGISTERS_reg[25][27]  ( .D(n3043), .CK(CLK), .Q(net310497), .QN(
        n17907) );
  DFF_X1 \REGISTERS_reg[25][26]  ( .D(n3042), .CK(CLK), .Q(net310496), .QN(
        n17906) );
  DFF_X1 \REGISTERS_reg[25][25]  ( .D(n3041), .CK(CLK), .Q(net310495), .QN(
        n17905) );
  DFF_X1 \REGISTERS_reg[25][24]  ( .D(n3040), .CK(CLK), .Q(net310494), .QN(
        n17904) );
  DFF_X1 \REGISTERS_reg[25][23]  ( .D(n3039), .CK(CLK), .Q(net310493), .QN(
        n17935) );
  DFF_X1 \REGISTERS_reg[25][22]  ( .D(n3038), .CK(CLK), .Q(net310492), .QN(
        n17934) );
  DFF_X1 \REGISTERS_reg[25][21]  ( .D(n3037), .CK(CLK), .Q(net310491), .QN(
        n17933) );
  DFF_X1 \REGISTERS_reg[25][20]  ( .D(n3036), .CK(CLK), .Q(net310490), .QN(
        n17932) );
  DFF_X1 \REGISTERS_reg[25][19]  ( .D(n3035), .CK(CLK), .Q(net310489), .QN(
        n17931) );
  DFF_X1 \REGISTERS_reg[25][18]  ( .D(n3034), .CK(CLK), .Q(net310488), .QN(
        n17930) );
  DFF_X1 \REGISTERS_reg[25][17]  ( .D(n3033), .CK(CLK), .Q(net310487), .QN(
        n17929) );
  DFF_X1 \REGISTERS_reg[25][16]  ( .D(n3032), .CK(CLK), .Q(net310486), .QN(
        n17928) );
  DFF_X1 \REGISTERS_reg[25][15]  ( .D(n3031), .CK(CLK), .Q(net310485), .QN(
        n17927) );
  DFF_X1 \REGISTERS_reg[25][14]  ( .D(n3030), .CK(CLK), .Q(net310484), .QN(
        n17926) );
  DFF_X1 \REGISTERS_reg[25][13]  ( .D(n3029), .CK(CLK), .Q(net310483), .QN(
        n17925) );
  DFF_X1 \REGISTERS_reg[25][12]  ( .D(n3028), .CK(CLK), .Q(net310482), .QN(
        n17924) );
  DFF_X1 \REGISTERS_reg[25][11]  ( .D(n3027), .CK(CLK), .Q(net310481), .QN(
        n17923) );
  DFF_X1 \REGISTERS_reg[25][10]  ( .D(n3026), .CK(CLK), .Q(net310480), .QN(
        n17922) );
  DFF_X1 \REGISTERS_reg[25][9]  ( .D(n3025), .CK(CLK), .Q(net310479), .QN(
        n17921) );
  DFF_X1 \REGISTERS_reg[25][8]  ( .D(n3024), .CK(CLK), .Q(net310478), .QN(
        n17920) );
  DFF_X1 \REGISTERS_reg[25][7]  ( .D(n3023), .CK(CLK), .Q(net310477), .QN(
        n17919) );
  DFF_X1 \REGISTERS_reg[25][6]  ( .D(n3022), .CK(CLK), .Q(net310476), .QN(
        n17918) );
  DFF_X1 \REGISTERS_reg[25][5]  ( .D(n3021), .CK(CLK), .Q(net310475), .QN(
        n17917) );
  DFF_X1 \REGISTERS_reg[25][4]  ( .D(n3020), .CK(CLK), .Q(net310474), .QN(
        n17916) );
  DFF_X1 \REGISTERS_reg[25][3]  ( .D(n3019), .CK(CLK), .Q(net310473), .QN(
        n17915) );
  DFF_X1 \REGISTERS_reg[25][2]  ( .D(n3018), .CK(CLK), .Q(net310472), .QN(
        n17913) );
  DFF_X1 \REGISTERS_reg[25][1]  ( .D(n3017), .CK(CLK), .Q(net310471), .QN(
        n17912) );
  DFF_X1 \REGISTERS_reg[25][0]  ( .D(n3016), .CK(CLK), .Q(net310470), .QN(
        n17914) );
  DFF_X1 \REGISTERS_reg[26][31]  ( .D(n3015), .CK(CLK), .QN(n17430) );
  DFF_X1 \REGISTERS_reg[26][30]  ( .D(n3014), .CK(CLK), .QN(n17429) );
  DFF_X1 \REGISTERS_reg[26][29]  ( .D(n3013), .CK(CLK), .QN(n17428) );
  DFF_X1 \REGISTERS_reg[26][28]  ( .D(n3012), .CK(CLK), .QN(n17427) );
  DFF_X1 \REGISTERS_reg[26][27]  ( .D(n3011), .CK(CLK), .QN(n17426) );
  DFF_X1 \REGISTERS_reg[26][26]  ( .D(n3010), .CK(CLK), .QN(n17425) );
  DFF_X1 \REGISTERS_reg[26][25]  ( .D(n3009), .CK(CLK), .QN(n17424) );
  DFF_X1 \REGISTERS_reg[26][24]  ( .D(n3008), .CK(CLK), .QN(n17423) );
  DFF_X1 \REGISTERS_reg[26][23]  ( .D(n3007), .CK(CLK), .QN(n17454) );
  DFF_X1 \REGISTERS_reg[26][22]  ( .D(n3006), .CK(CLK), .QN(n17453) );
  DFF_X1 \REGISTERS_reg[26][21]  ( .D(n3005), .CK(CLK), .QN(n17452) );
  DFF_X1 \REGISTERS_reg[26][20]  ( .D(n3004), .CK(CLK), .QN(n17451) );
  DFF_X1 \REGISTERS_reg[26][19]  ( .D(n3003), .CK(CLK), .QN(n17450) );
  DFF_X1 \REGISTERS_reg[26][18]  ( .D(n3002), .CK(CLK), .QN(n17449) );
  DFF_X1 \REGISTERS_reg[26][17]  ( .D(n3001), .CK(CLK), .QN(n17448) );
  DFF_X1 \REGISTERS_reg[26][16]  ( .D(n3000), .CK(CLK), .QN(n17447) );
  DFF_X1 \REGISTERS_reg[26][15]  ( .D(n2999), .CK(CLK), .QN(n17446) );
  DFF_X1 \REGISTERS_reg[26][14]  ( .D(n2998), .CK(CLK), .QN(n17445) );
  DFF_X1 \REGISTERS_reg[26][13]  ( .D(n2997), .CK(CLK), .QN(n17444) );
  DFF_X1 \REGISTERS_reg[26][12]  ( .D(n2996), .CK(CLK), .QN(n17443) );
  DFF_X1 \REGISTERS_reg[26][11]  ( .D(n2995), .CK(CLK), .QN(n17442) );
  DFF_X1 \REGISTERS_reg[26][10]  ( .D(n2994), .CK(CLK), .QN(n17441) );
  DFF_X1 \REGISTERS_reg[26][9]  ( .D(n2993), .CK(CLK), .QN(n17440) );
  DFF_X1 \REGISTERS_reg[26][8]  ( .D(n2992), .CK(CLK), .QN(n17439) );
  DFF_X1 \REGISTERS_reg[26][7]  ( .D(n2991), .CK(CLK), .QN(n17438) );
  DFF_X1 \REGISTERS_reg[26][6]  ( .D(n2990), .CK(CLK), .QN(n17437) );
  DFF_X1 \REGISTERS_reg[26][5]  ( .D(n2989), .CK(CLK), .QN(n17436) );
  DFF_X1 \REGISTERS_reg[26][4]  ( .D(n2988), .CK(CLK), .QN(n17435) );
  DFF_X1 \REGISTERS_reg[26][3]  ( .D(n2987), .CK(CLK), .QN(n17434) );
  DFF_X1 \REGISTERS_reg[26][2]  ( .D(n2986), .CK(CLK), .QN(n17432) );
  DFF_X1 \REGISTERS_reg[26][1]  ( .D(n2985), .CK(CLK), .QN(n17433) );
  DFF_X1 \REGISTERS_reg[26][0]  ( .D(n2984), .CK(CLK), .QN(n17431) );
  DFF_X1 \REGISTERS_reg[27][31]  ( .D(n2983), .CK(CLK), .QN(n17668) );
  DFF_X1 \REGISTERS_reg[27][30]  ( .D(n2982), .CK(CLK), .QN(n17667) );
  DFF_X1 \REGISTERS_reg[27][29]  ( .D(n2981), .CK(CLK), .QN(n17666) );
  DFF_X1 \REGISTERS_reg[27][28]  ( .D(n2980), .CK(CLK), .QN(n17665) );
  DFF_X1 \REGISTERS_reg[27][27]  ( .D(n2979), .CK(CLK), .QN(n17664) );
  DFF_X1 \REGISTERS_reg[27][26]  ( .D(n2978), .CK(CLK), .QN(n17663) );
  DFF_X1 \REGISTERS_reg[27][25]  ( .D(n2977), .CK(CLK), .QN(n17662) );
  DFF_X1 \REGISTERS_reg[27][24]  ( .D(n2976), .CK(CLK), .QN(n17661) );
  DFF_X1 \REGISTERS_reg[27][23]  ( .D(n2975), .CK(CLK), .QN(n17660) );
  DFF_X1 \REGISTERS_reg[27][22]  ( .D(n2974), .CK(CLK), .QN(n17659) );
  DFF_X1 \REGISTERS_reg[27][21]  ( .D(n2973), .CK(CLK), .QN(n17658) );
  DFF_X1 \REGISTERS_reg[27][20]  ( .D(n2972), .CK(CLK), .QN(n17657) );
  DFF_X1 \REGISTERS_reg[27][19]  ( .D(n2971), .CK(CLK), .QN(n17656) );
  DFF_X1 \REGISTERS_reg[27][18]  ( .D(n2970), .CK(CLK), .QN(n17655) );
  DFF_X1 \REGISTERS_reg[27][17]  ( .D(n2969), .CK(CLK), .QN(n17654) );
  DFF_X1 \REGISTERS_reg[27][16]  ( .D(n2968), .CK(CLK), .QN(n17653) );
  DFF_X1 \REGISTERS_reg[27][15]  ( .D(n2967), .CK(CLK), .QN(n17652) );
  DFF_X1 \REGISTERS_reg[27][14]  ( .D(n2966), .CK(CLK), .QN(n17651) );
  DFF_X1 \REGISTERS_reg[27][13]  ( .D(n2965), .CK(CLK), .QN(n17650) );
  DFF_X1 \REGISTERS_reg[27][12]  ( .D(n2964), .CK(CLK), .QN(n17649) );
  DFF_X1 \REGISTERS_reg[27][11]  ( .D(n2963), .CK(CLK), .QN(n17648) );
  DFF_X1 \REGISTERS_reg[27][10]  ( .D(n2962), .CK(CLK), .QN(n17647) );
  DFF_X1 \REGISTERS_reg[27][9]  ( .D(n2961), .CK(CLK), .QN(n17646) );
  DFF_X1 \REGISTERS_reg[27][8]  ( .D(n2960), .CK(CLK), .QN(n17645) );
  DFF_X1 \REGISTERS_reg[27][7]  ( .D(n2959), .CK(CLK), .QN(n17644) );
  DFF_X1 \REGISTERS_reg[27][6]  ( .D(n2958), .CK(CLK), .QN(n17643) );
  DFF_X1 \REGISTERS_reg[27][5]  ( .D(n2957), .CK(CLK), .QN(n17642) );
  DFF_X1 \REGISTERS_reg[27][4]  ( .D(n2956), .CK(CLK), .QN(n17641) );
  DFF_X1 \REGISTERS_reg[27][3]  ( .D(n2955), .CK(CLK), .QN(n17640) );
  DFF_X1 \REGISTERS_reg[27][2]  ( .D(n2954), .CK(CLK), .QN(n17678) );
  DFF_X1 \REGISTERS_reg[27][1]  ( .D(n2953), .CK(CLK), .QN(n17639) );
  DFF_X1 \REGISTERS_reg[27][0]  ( .D(n2952), .CK(CLK), .QN(n17638) );
  DFF_X1 \REGISTERS_reg[28][31]  ( .D(n2951), .CK(CLK), .QN(n17526) );
  DFF_X1 \REGISTERS_reg[28][30]  ( .D(n2950), .CK(CLK), .QN(n17525) );
  DFF_X1 \REGISTERS_reg[28][29]  ( .D(n2949), .CK(CLK), .QN(n17524) );
  DFF_X1 \REGISTERS_reg[28][28]  ( .D(n2948), .CK(CLK), .QN(n17523) );
  DFF_X1 \REGISTERS_reg[28][27]  ( .D(n2947), .CK(CLK), .QN(n17522) );
  DFF_X1 \REGISTERS_reg[28][26]  ( .D(n2946), .CK(CLK), .QN(n17521) );
  DFF_X1 \REGISTERS_reg[28][25]  ( .D(n2945), .CK(CLK), .QN(n17520) );
  DFF_X1 \REGISTERS_reg[28][24]  ( .D(n2944), .CK(CLK), .QN(n17519) );
  DFF_X1 \REGISTERS_reg[28][23]  ( .D(n2943), .CK(CLK), .QN(n17561) );
  DFF_X1 \REGISTERS_reg[28][22]  ( .D(n2942), .CK(CLK), .QN(n17560) );
  DFF_X1 \REGISTERS_reg[28][21]  ( .D(n2941), .CK(CLK), .QN(n17559) );
  DFF_X1 \REGISTERS_reg[28][20]  ( .D(n2940), .CK(CLK), .QN(n17558) );
  DFF_X1 \REGISTERS_reg[28][19]  ( .D(n2939), .CK(CLK), .QN(n17557) );
  DFF_X1 \REGISTERS_reg[28][18]  ( .D(n2938), .CK(CLK), .QN(n17556) );
  DFF_X1 \REGISTERS_reg[28][17]  ( .D(n2937), .CK(CLK), .QN(n17555) );
  DFF_X1 \REGISTERS_reg[28][16]  ( .D(n2936), .CK(CLK), .QN(n17554) );
  DFF_X1 \REGISTERS_reg[28][15]  ( .D(n2935), .CK(CLK), .QN(n17553) );
  DFF_X1 \REGISTERS_reg[28][14]  ( .D(n2934), .CK(CLK), .QN(n17552) );
  DFF_X1 \REGISTERS_reg[28][13]  ( .D(n2933), .CK(CLK), .QN(n17551) );
  DFF_X1 \REGISTERS_reg[28][12]  ( .D(n2932), .CK(CLK), .QN(n17550) );
  DFF_X1 \REGISTERS_reg[28][11]  ( .D(n2931), .CK(CLK), .QN(n17549) );
  DFF_X1 \REGISTERS_reg[28][10]  ( .D(n2930), .CK(CLK), .QN(n17548) );
  DFF_X1 \REGISTERS_reg[28][9]  ( .D(n2929), .CK(CLK), .QN(n17547) );
  DFF_X1 \REGISTERS_reg[28][8]  ( .D(n2928), .CK(CLK), .QN(n17546) );
  DFF_X1 \REGISTERS_reg[28][7]  ( .D(n2927), .CK(CLK), .QN(n17545) );
  DFF_X1 \REGISTERS_reg[28][6]  ( .D(n2926), .CK(CLK), .QN(n17544) );
  DFF_X1 \REGISTERS_reg[28][5]  ( .D(n2925), .CK(CLK), .QN(n17543) );
  DFF_X1 \REGISTERS_reg[28][4]  ( .D(n2924), .CK(CLK), .QN(n17542) );
  DFF_X1 \REGISTERS_reg[28][3]  ( .D(n2923), .CK(CLK), .QN(n17541) );
  DFF_X1 \REGISTERS_reg[28][2]  ( .D(n2922), .CK(CLK), .QN(n17540) );
  DFF_X1 \REGISTERS_reg[28][1]  ( .D(n2921), .CK(CLK), .QN(n17536) );
  DFF_X1 \REGISTERS_reg[28][0]  ( .D(n2920), .CK(CLK), .QN(n17535) );
  DFF_X1 \REGISTERS_reg[29][31]  ( .D(n2919), .CK(CLK), .QN(n17613) );
  DFF_X1 \REGISTERS_reg[29][30]  ( .D(n2918), .CK(CLK), .QN(n17612) );
  DFF_X1 \REGISTERS_reg[29][29]  ( .D(n2917), .CK(CLK), .QN(n17611) );
  DFF_X1 \REGISTERS_reg[29][28]  ( .D(n2916), .CK(CLK), .QN(n17610) );
  DFF_X1 \REGISTERS_reg[29][27]  ( .D(n2915), .CK(CLK), .QN(n17609) );
  DFF_X1 \REGISTERS_reg[29][26]  ( .D(n2914), .CK(CLK), .QN(n17608) );
  DFF_X1 \REGISTERS_reg[29][25]  ( .D(n2913), .CK(CLK), .QN(n17607) );
  DFF_X1 \REGISTERS_reg[29][24]  ( .D(n2912), .CK(CLK), .QN(n17606) );
  DFF_X1 \REGISTERS_reg[29][23]  ( .D(n2911), .CK(CLK), .QN(n17605) );
  DFF_X1 \REGISTERS_reg[29][22]  ( .D(n2910), .CK(CLK), .QN(n17604) );
  DFF_X1 \REGISTERS_reg[29][21]  ( .D(n2909), .CK(CLK), .QN(n17603) );
  DFF_X1 \REGISTERS_reg[29][20]  ( .D(n2908), .CK(CLK), .QN(n17602) );
  DFF_X1 \REGISTERS_reg[29][19]  ( .D(n2907), .CK(CLK), .QN(n17601) );
  DFF_X1 \REGISTERS_reg[29][18]  ( .D(n2906), .CK(CLK), .QN(n17600) );
  DFF_X1 \REGISTERS_reg[29][17]  ( .D(n2905), .CK(CLK), .QN(n17599) );
  DFF_X1 \REGISTERS_reg[29][16]  ( .D(n2904), .CK(CLK), .QN(n17598) );
  DFF_X1 \REGISTERS_reg[29][15]  ( .D(n2903), .CK(CLK), .QN(n17597) );
  DFF_X1 \REGISTERS_reg[29][14]  ( .D(n2902), .CK(CLK), .QN(n17596) );
  DFF_X1 \REGISTERS_reg[29][13]  ( .D(n2901), .CK(CLK), .QN(n17595) );
  DFF_X1 \REGISTERS_reg[29][12]  ( .D(n2900), .CK(CLK), .QN(n17594) );
  DFF_X1 \REGISTERS_reg[29][11]  ( .D(n2899), .CK(CLK), .QN(n17593) );
  DFF_X1 \REGISTERS_reg[29][10]  ( .D(n2898), .CK(CLK), .QN(n17592) );
  DFF_X1 \REGISTERS_reg[29][9]  ( .D(n2897), .CK(CLK), .QN(n17591) );
  DFF_X1 \REGISTERS_reg[29][8]  ( .D(n2896), .CK(CLK), .QN(n17590) );
  DFF_X1 \REGISTERS_reg[29][7]  ( .D(n2895), .CK(CLK), .QN(n17589) );
  DFF_X1 \REGISTERS_reg[29][6]  ( .D(n2894), .CK(CLK), .QN(n17588) );
  DFF_X1 \REGISTERS_reg[29][5]  ( .D(n2893), .CK(CLK), .QN(n17587) );
  DFF_X1 \REGISTERS_reg[29][4]  ( .D(n2892), .CK(CLK), .QN(n17586) );
  DFF_X1 \REGISTERS_reg[29][3]  ( .D(n2891), .CK(CLK), .QN(n17585) );
  DFF_X1 \REGISTERS_reg[29][2]  ( .D(n2890), .CK(CLK), .QN(n17584) );
  DFF_X1 \REGISTERS_reg[29][1]  ( .D(n2889), .CK(CLK), .QN(n17677) );
  DFF_X1 \REGISTERS_reg[29][0]  ( .D(n2888), .CK(CLK), .QN(n17583) );
  DFF_X1 \REGISTERS_reg[30][31]  ( .D(n2887), .CK(CLK), .QN(n17494) );
  DFF_X1 \REGISTERS_reg[30][30]  ( .D(n2886), .CK(CLK), .QN(n17493) );
  DFF_X1 \REGISTERS_reg[30][29]  ( .D(n2885), .CK(CLK), .QN(n17492) );
  DFF_X1 \REGISTERS_reg[30][28]  ( .D(n2884), .CK(CLK), .QN(n17491) );
  DFF_X1 \REGISTERS_reg[30][27]  ( .D(n2883), .CK(CLK), .QN(n17490) );
  DFF_X1 \REGISTERS_reg[30][26]  ( .D(n2882), .CK(CLK), .QN(n17489) );
  DFF_X1 \REGISTERS_reg[30][25]  ( .D(n2881), .CK(CLK), .QN(n17488) );
  DFF_X1 \REGISTERS_reg[30][24]  ( .D(n2880), .CK(CLK), .QN(n17487) );
  DFF_X1 \REGISTERS_reg[30][23]  ( .D(n2879), .CK(CLK), .QN(n17517) );
  DFF_X1 \REGISTERS_reg[30][22]  ( .D(n2878), .CK(CLK), .QN(n17516) );
  DFF_X1 \REGISTERS_reg[30][21]  ( .D(n2877), .CK(CLK), .QN(n17515) );
  DFF_X1 \REGISTERS_reg[30][20]  ( .D(n2876), .CK(CLK), .QN(n17514) );
  DFF_X1 \REGISTERS_reg[30][19]  ( .D(n2875), .CK(CLK), .QN(n17513) );
  DFF_X1 \REGISTERS_reg[30][18]  ( .D(n2874), .CK(CLK), .QN(n17512) );
  DFF_X1 \REGISTERS_reg[30][17]  ( .D(n2873), .CK(CLK), .QN(n17511) );
  DFF_X1 \REGISTERS_reg[30][16]  ( .D(n2872), .CK(CLK), .QN(n17510) );
  DFF_X1 \REGISTERS_reg[30][15]  ( .D(n2871), .CK(CLK), .QN(n17509) );
  DFF_X1 \REGISTERS_reg[30][14]  ( .D(n2870), .CK(CLK), .QN(n17508) );
  DFF_X1 \REGISTERS_reg[30][13]  ( .D(n2869), .CK(CLK), .QN(n17507) );
  DFF_X1 \REGISTERS_reg[30][12]  ( .D(n2868), .CK(CLK), .QN(n17506) );
  DFF_X1 \REGISTERS_reg[30][11]  ( .D(n2867), .CK(CLK), .QN(n17505) );
  DFF_X1 \REGISTERS_reg[30][10]  ( .D(n2866), .CK(CLK), .QN(n17504) );
  DFF_X1 \REGISTERS_reg[30][9]  ( .D(n2865), .CK(CLK), .QN(n17503) );
  DFF_X1 \REGISTERS_reg[30][8]  ( .D(n2864), .CK(CLK), .QN(n17502) );
  DFF_X1 \REGISTERS_reg[30][7]  ( .D(n2863), .CK(CLK), .QN(n17501) );
  DFF_X1 \REGISTERS_reg[30][6]  ( .D(n2862), .CK(CLK), .QN(n17500) );
  DFF_X1 \REGISTERS_reg[30][5]  ( .D(n2861), .CK(CLK), .QN(n17499) );
  DFF_X1 \REGISTERS_reg[30][4]  ( .D(n2860), .CK(CLK), .QN(n17498) );
  DFF_X1 \REGISTERS_reg[30][3]  ( .D(n2859), .CK(CLK), .QN(n17497) );
  DFF_X1 \REGISTERS_reg[30][2]  ( .D(n2858), .CK(CLK), .QN(n17496) );
  DFF_X1 \REGISTERS_reg[30][1]  ( .D(n2857), .CK(CLK), .QN(n17495) );
  DFF_X1 \REGISTERS_reg[30][0]  ( .D(n2856), .CK(CLK), .QN(n17518) );
  DFF_X1 \REGISTERS_reg[31][31]  ( .D(n2855), .CK(CLK), .Q(net591562), .QN(
        n18320) );
  DFF_X1 \OUT1_reg[31]  ( .D(n2854), .CK(CLK), .Q(OUT1[31]) );
  DFF_X1 \REGISTERS_reg[31][30]  ( .D(n2853), .CK(CLK), .Q(net591561), .QN(
        n18326) );
  DFF_X1 \OUT1_reg[30]  ( .D(n2852), .CK(CLK), .Q(OUT1[30]) );
  DFF_X1 \REGISTERS_reg[31][29]  ( .D(n2851), .CK(CLK), .Q(net591560), .QN(
        n18325) );
  DFF_X1 \OUT1_reg[29]  ( .D(n2850), .CK(CLK), .Q(OUT1[29]) );
  DFF_X1 \REGISTERS_reg[31][28]  ( .D(n2849), .CK(CLK), .Q(net591559), .QN(
        n18324) );
  DFF_X1 \OUT1_reg[28]  ( .D(n2848), .CK(CLK), .Q(OUT1[28]) );
  DFF_X1 \REGISTERS_reg[31][27]  ( .D(n2847), .CK(CLK), .Q(net591558), .QN(
        n18323) );
  DFF_X1 \OUT1_reg[27]  ( .D(n2846), .CK(CLK), .Q(OUT1[27]) );
  DFF_X1 \REGISTERS_reg[31][26]  ( .D(n2845), .CK(CLK), .Q(net591557), .QN(
        n18322) );
  DFF_X1 \OUT1_reg[26]  ( .D(n2844), .CK(CLK), .Q(OUT1[26]) );
  DFF_X1 \REGISTERS_reg[31][25]  ( .D(n2843), .CK(CLK), .Q(net591556), .QN(
        n18321) );
  DFF_X1 \OUT1_reg[25]  ( .D(n2842), .CK(CLK), .Q(OUT1[25]) );
  DFF_X1 \REGISTERS_reg[31][24]  ( .D(n2841), .CK(CLK), .Q(net591555), .QN(
        n18339) );
  DFF_X1 \OUT1_reg[24]  ( .D(n2840), .CK(CLK), .Q(OUT1[24]) );
  DFF_X1 \REGISTERS_reg[31][23]  ( .D(n2839), .CK(CLK), .Q(net591554), .QN(
        n18338) );
  DFF_X1 \OUT1_reg[23]  ( .D(n2838), .CK(CLK), .Q(OUT1[23]) );
  DFF_X1 \REGISTERS_reg[31][22]  ( .D(n2837), .CK(CLK), .Q(net591553), .QN(
        n18337) );
  DFF_X1 \OUT1_reg[22]  ( .D(n2836), .CK(CLK), .Q(OUT1[22]) );
  DFF_X1 \REGISTERS_reg[31][21]  ( .D(n2835), .CK(CLK), .Q(net591552), .QN(
        n18336) );
  DFF_X1 \OUT1_reg[21]  ( .D(n2834), .CK(CLK), .Q(OUT1[21]) );
  DFF_X1 \REGISTERS_reg[31][20]  ( .D(n2833), .CK(CLK), .Q(net591551), .QN(
        n18335) );
  DFF_X1 \OUT1_reg[20]  ( .D(n2832), .CK(CLK), .Q(OUT1[20]) );
  DFF_X1 \REGISTERS_reg[31][19]  ( .D(n2831), .CK(CLK), .Q(net591550), .QN(
        n18334) );
  DFF_X1 \OUT1_reg[19]  ( .D(n2830), .CK(CLK), .Q(OUT1[19]) );
  DFF_X1 \REGISTERS_reg[31][18]  ( .D(n2829), .CK(CLK), .Q(net591549), .QN(
        n18333) );
  DFF_X1 \OUT1_reg[18]  ( .D(n2828), .CK(CLK), .Q(OUT1[18]) );
  DFF_X1 \REGISTERS_reg[31][17]  ( .D(n2827), .CK(CLK), .Q(net591548), .QN(
        n18332) );
  DFF_X1 \OUT1_reg[17]  ( .D(n2826), .CK(CLK), .Q(OUT1[17]) );
  DFF_X1 \REGISTERS_reg[31][16]  ( .D(n2825), .CK(CLK), .Q(net591547), .QN(
        n18331) );
  DFF_X1 \OUT1_reg[16]  ( .D(n2824), .CK(CLK), .Q(OUT1[16]) );
  DFF_X1 \REGISTERS_reg[31][15]  ( .D(n2823), .CK(CLK), .Q(net591546), .QN(
        n18330) );
  DFF_X1 \OUT1_reg[15]  ( .D(n2822), .CK(CLK), .Q(OUT1[15]) );
  DFF_X1 \REGISTERS_reg[31][14]  ( .D(n2821), .CK(CLK), .Q(net591545), .QN(
        n18329) );
  DFF_X1 \OUT1_reg[14]  ( .D(n2820), .CK(CLK), .Q(OUT1[14]) );
  DFF_X1 \REGISTERS_reg[31][13]  ( .D(n2819), .CK(CLK), .Q(net591544), .QN(
        n18328) );
  DFF_X1 \OUT1_reg[13]  ( .D(n2818), .CK(CLK), .Q(OUT1[13]) );
  DFF_X1 \REGISTERS_reg[31][12]  ( .D(n2817), .CK(CLK), .Q(net591543), .QN(
        n18327) );
  DFF_X1 \OUT1_reg[12]  ( .D(n2816), .CK(CLK), .Q(OUT1[12]) );
  DFF_X1 \REGISTERS_reg[31][11]  ( .D(n2815), .CK(CLK), .Q(net591542), .QN(
        n18346) );
  DFF_X1 \OUT1_reg[11]  ( .D(n2814), .CK(CLK), .Q(OUT1[11]) );
  DFF_X1 \REGISTERS_reg[31][10]  ( .D(n2813), .CK(CLK), .Q(net591541), .QN(
        n18345) );
  DFF_X1 \OUT1_reg[10]  ( .D(n2812), .CK(CLK), .Q(OUT1[10]) );
  DFF_X1 \REGISTERS_reg[31][9]  ( .D(n2811), .CK(CLK), .Q(net591540), .QN(
        n18344) );
  DFF_X1 \OUT1_reg[9]  ( .D(n2810), .CK(CLK), .Q(OUT1[9]) );
  DFF_X1 \REGISTERS_reg[31][8]  ( .D(n2809), .CK(CLK), .Q(net591539), .QN(
        n18343) );
  DFF_X1 \OUT1_reg[8]  ( .D(n2808), .CK(CLK), .Q(OUT1[8]) );
  DFF_X1 \REGISTERS_reg[31][7]  ( .D(n2807), .CK(CLK), .Q(net591538), .QN(
        n18342) );
  DFF_X1 \OUT1_reg[7]  ( .D(n2806), .CK(CLK), .Q(OUT1[7]) );
  DFF_X1 \REGISTERS_reg[31][6]  ( .D(n2805), .CK(CLK), .Q(net591537), .QN(
        n18341) );
  DFF_X1 \OUT1_reg[6]  ( .D(n2804), .CK(CLK), .Q(OUT1[6]) );
  DFF_X1 \REGISTERS_reg[31][5]  ( .D(n2803), .CK(CLK), .Q(net591536), .QN(
        n18340) );
  DFF_X1 \OUT1_reg[5]  ( .D(n2802), .CK(CLK), .Q(OUT1[5]) );
  DFF_X1 \REGISTERS_reg[31][4]  ( .D(n2801), .CK(CLK), .Q(net591535), .QN(
        n18351) );
  DFF_X1 \OUT1_reg[4]  ( .D(n2800), .CK(CLK), .Q(OUT1[4]) );
  DFF_X1 \REGISTERS_reg[31][3]  ( .D(n2799), .CK(CLK), .Q(net591534), .QN(
        n18350) );
  DFF_X1 \OUT1_reg[3]  ( .D(n2798), .CK(CLK), .Q(OUT1[3]) );
  DFF_X1 \REGISTERS_reg[31][2]  ( .D(n2797), .CK(CLK), .Q(net591533), .QN(
        n18349) );
  DFF_X1 \OUT1_reg[2]  ( .D(n2796), .CK(CLK), .Q(OUT1[2]) );
  DFF_X1 \REGISTERS_reg[31][1]  ( .D(n2795), .CK(CLK), .Q(net591532), .QN(
        n18348) );
  DFF_X1 \OUT1_reg[1]  ( .D(n2794), .CK(CLK), .Q(OUT1[1]) );
  DFF_X1 \REGISTERS_reg[31][0]  ( .D(n2793), .CK(CLK), .Q(net591531), .QN(
        n18347) );
  DFF_X1 \OUT1_reg[0]  ( .D(n2792), .CK(CLK), .Q(OUT1[0]) );
  DFF_X1 \OUT2_reg[31]  ( .D(n2791), .CK(CLK), .Q(OUT2[31]) );
  DFF_X1 \OUT2_reg[30]  ( .D(n2790), .CK(CLK), .Q(OUT2[30]) );
  DFF_X1 \OUT2_reg[29]  ( .D(n2789), .CK(CLK), .Q(OUT2[29]) );
  DFF_X1 \OUT2_reg[28]  ( .D(n2788), .CK(CLK), .Q(OUT2[28]) );
  DFF_X1 \OUT2_reg[27]  ( .D(n2787), .CK(CLK), .Q(OUT2[27]) );
  DFF_X1 \OUT2_reg[26]  ( .D(n2786), .CK(CLK), .Q(OUT2[26]) );
  DFF_X1 \OUT2_reg[25]  ( .D(n2785), .CK(CLK), .Q(OUT2[25]) );
  DFF_X1 \OUT2_reg[24]  ( .D(n2784), .CK(CLK), .Q(OUT2[24]) );
  DFF_X1 \OUT2_reg[23]  ( .D(n2783), .CK(CLK), .Q(OUT2[23]) );
  DFF_X1 \OUT2_reg[22]  ( .D(n2782), .CK(CLK), .Q(OUT2[22]) );
  DFF_X1 \OUT2_reg[21]  ( .D(n2781), .CK(CLK), .Q(OUT2[21]) );
  DFF_X1 \OUT2_reg[20]  ( .D(n2780), .CK(CLK), .Q(OUT2[20]) );
  DFF_X1 \OUT2_reg[19]  ( .D(n2779), .CK(CLK), .Q(OUT2[19]) );
  DFF_X1 \OUT2_reg[18]  ( .D(n2778), .CK(CLK), .Q(OUT2[18]) );
  DFF_X1 \OUT2_reg[17]  ( .D(n2777), .CK(CLK), .Q(OUT2[17]) );
  DFF_X1 \OUT2_reg[16]  ( .D(n2776), .CK(CLK), .Q(OUT2[16]) );
  DFF_X1 \OUT2_reg[15]  ( .D(n2775), .CK(CLK), .Q(OUT2[15]) );
  DFF_X1 \OUT2_reg[14]  ( .D(n2774), .CK(CLK), .Q(OUT2[14]) );
  DFF_X1 \OUT2_reg[13]  ( .D(n2773), .CK(CLK), .Q(OUT2[13]) );
  DFF_X1 \OUT2_reg[12]  ( .D(n2772), .CK(CLK), .Q(OUT2[12]) );
  DFF_X1 \OUT2_reg[11]  ( .D(n2771), .CK(CLK), .Q(OUT2[11]) );
  DFF_X1 \OUT2_reg[10]  ( .D(n2770), .CK(CLK), .Q(OUT2[10]) );
  DFF_X1 \OUT2_reg[9]  ( .D(n2769), .CK(CLK), .Q(OUT2[9]) );
  DFF_X1 \OUT2_reg[8]  ( .D(n2768), .CK(CLK), .Q(OUT2[8]) );
  DFF_X1 \OUT2_reg[7]  ( .D(n2767), .CK(CLK), .Q(OUT2[7]) );
  DFF_X1 \OUT2_reg[6]  ( .D(n2766), .CK(CLK), .Q(OUT2[6]) );
  DFF_X1 \OUT2_reg[5]  ( .D(n2765), .CK(CLK), .Q(OUT2[5]) );
  DFF_X1 \OUT2_reg[4]  ( .D(n2764), .CK(CLK), .Q(OUT2[4]) );
  DFF_X1 \OUT2_reg[3]  ( .D(n2763), .CK(CLK), .Q(OUT2[3]) );
  DFF_X1 \OUT2_reg[2]  ( .D(n2762), .CK(CLK), .Q(OUT2[2]) );
  DFF_X1 \OUT2_reg[1]  ( .D(n2761), .CK(CLK), .Q(OUT2[1]) );
  DFF_X1 \OUT2_reg[0]  ( .D(n2760), .CK(CLK), .Q(OUT2[0]) );
  NAND3_X1 U3477 ( .A1(n1248), .A2(n1249), .A3(n1250), .ZN(n1138) );
  NAND3_X1 U3478 ( .A1(n1250), .A2(n1249), .A3(ADD_WR[2]), .ZN(n1286) );
  NAND3_X1 U3479 ( .A1(n1250), .A2(n1248), .A3(ADD_WR[3]), .ZN(n1424) );
  NAND3_X1 U3480 ( .A1(ADD_WR[2]), .A2(n1250), .A3(ADD_WR[3]), .ZN(n1561) );
  NAND3_X1 U3481 ( .A1(n1248), .A2(n1249), .A3(n1803), .ZN(n1700) );
  NAND3_X1 U3482 ( .A1(ADD_WR[2]), .A2(n1249), .A3(n1803), .ZN(n1838) );
  NAND3_X1 U3483 ( .A1(ADD_WR[3]), .A2(n1248), .A3(n1803), .ZN(n1975) );
  NAND3_X1 U3484 ( .A1(ADD_WR[3]), .A2(ADD_WR[2]), .A3(n1803), .ZN(n2112) );
  NOR3_X1 U3 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .A3(n18441), .ZN(n4543) );
  NOR3_X1 U4 ( .A1(n18441), .A2(ADD_RD2[1]), .A3(n4553), .ZN(n4532) );
  NOR3_X1 U5 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .A3(n18539), .ZN(n3906) );
  NOR3_X1 U6 ( .A1(n18538), .A2(ADD_RD1[2]), .A3(n3925), .ZN(n3917) );
  NOR2_X2 U7 ( .A1(DATAIN[4]), .A2(n18994), .ZN(n1694) );
  NOR2_X2 U8 ( .A1(DATAIN[3]), .A2(n18994), .ZN(n1419) );
  NOR2_X2 U9 ( .A1(DATAIN[2]), .A2(n18994), .ZN(n1282) );
  NOR2_X2 U10 ( .A1(DATAIN[1]), .A2(n18995), .ZN(n1209) );
  NOR2_X2 U11 ( .A1(DATAIN[0]), .A2(n18995), .ZN(n1174) );
  NAND2_X1 U12 ( .A1(DATAIN[0]), .A2(n18997), .ZN(n1136) );
  NAND2_X1 U13 ( .A1(DATAIN[1]), .A2(n18997), .ZN(n1134) );
  NAND2_X1 U14 ( .A1(DATAIN[2]), .A2(n18997), .ZN(n1132) );
  NAND2_X1 U15 ( .A1(DATAIN[3]), .A2(n18997), .ZN(n1130) );
  NAND2_X1 U16 ( .A1(DATAIN[4]), .A2(n18997), .ZN(n1128) );
  AND3_X1 U17 ( .A1(ENABLE), .A2(n18998), .A3(RD2), .ZN(n17839) );
  INV_X1 U18 ( .A(n18734), .ZN(n18725) );
  BUF_X1 U19 ( .A(n3963), .Z(n18401) );
  BUF_X1 U20 ( .A(n3967), .Z(n18389) );
  BUF_X1 U21 ( .A(n3963), .Z(n18402) );
  BUF_X1 U22 ( .A(n3967), .Z(n18390) );
  BUF_X1 U23 ( .A(n3975), .Z(n18368) );
  BUF_X1 U24 ( .A(n3980), .Z(n18356) );
  BUF_X1 U25 ( .A(n3975), .Z(n18369) );
  BUF_X1 U26 ( .A(n3980), .Z(n18357) );
  BUF_X1 U27 ( .A(n3976), .Z(n18365) );
  BUF_X1 U28 ( .A(n3976), .Z(n18366) );
  BUF_X1 U29 ( .A(n3964), .Z(n18398) );
  BUF_X1 U30 ( .A(n3981), .Z(n18353) );
  BUF_X1 U31 ( .A(n3964), .Z(n18399) );
  BUF_X1 U32 ( .A(n3981), .Z(n18354) );
  BUF_X1 U33 ( .A(n3940), .Z(n18445) );
  BUF_X1 U34 ( .A(n3940), .Z(n18446) );
  BUF_X1 U35 ( .A(n3945), .Z(n18434) );
  BUF_X1 U36 ( .A(n3945), .Z(n18435) );
  BUF_X1 U37 ( .A(n3977), .Z(n18362) );
  BUF_X1 U38 ( .A(n3977), .Z(n18363) );
  BUF_X1 U39 ( .A(n3957), .Z(n18407) );
  BUF_X1 U40 ( .A(n3942), .Z(n18442) );
  BUF_X1 U41 ( .A(n3957), .Z(n18408) );
  BUF_X1 U42 ( .A(n3942), .Z(n18443) );
  BUF_X1 U43 ( .A(n3978), .Z(n18359) );
  BUF_X1 U44 ( .A(n3978), .Z(n18360) );
  BUF_X1 U45 ( .A(n3949), .Z(n18425) );
  BUF_X1 U46 ( .A(n3949), .Z(n18426) );
  BUF_X1 U47 ( .A(n3963), .Z(n18403) );
  BUF_X1 U48 ( .A(n3967), .Z(n18391) );
  BUF_X1 U49 ( .A(n3975), .Z(n18370) );
  BUF_X1 U50 ( .A(n3980), .Z(n18358) );
  BUF_X1 U51 ( .A(n3969), .Z(n18383) );
  BUF_X1 U52 ( .A(n3969), .Z(n18384) );
  BUF_X1 U53 ( .A(n3976), .Z(n18367) );
  BUF_X1 U54 ( .A(n3964), .Z(n18400) );
  BUF_X1 U55 ( .A(n3981), .Z(n18355) );
  BUF_X1 U56 ( .A(n3958), .Z(n18405) );
  BUF_X1 U57 ( .A(n3958), .Z(n18404) );
  BUF_X1 U58 ( .A(n3940), .Z(n18447) );
  BUF_X1 U59 ( .A(n3945), .Z(n18436) );
  BUF_X1 U60 ( .A(n3977), .Z(n18364) );
  BUF_X1 U61 ( .A(n3957), .Z(n18409) );
  BUF_X1 U62 ( .A(n3942), .Z(n18444) );
  BUF_X1 U63 ( .A(n3978), .Z(n18361) );
  BUF_X1 U64 ( .A(n3949), .Z(n18427) );
  BUF_X1 U65 ( .A(n3969), .Z(n18385) );
  BUF_X1 U66 ( .A(n3958), .Z(n18406) );
  INV_X1 U67 ( .A(n18596), .ZN(n18586) );
  INV_X1 U68 ( .A(n18596), .ZN(n18587) );
  INV_X1 U69 ( .A(n18621), .ZN(n18612) );
  INV_X1 U70 ( .A(n18632), .ZN(n18623) );
  INV_X1 U71 ( .A(n18643), .ZN(n18634) );
  INV_X1 U72 ( .A(n18668), .ZN(n18659) );
  INV_X1 U73 ( .A(n18679), .ZN(n18670) );
  INV_X1 U74 ( .A(n18690), .ZN(n18681) );
  INV_X1 U75 ( .A(n18701), .ZN(n18692) );
  INV_X1 U76 ( .A(n18712), .ZN(n18703) );
  INV_X1 U77 ( .A(n18723), .ZN(n18714) );
  INV_X1 U78 ( .A(n18759), .ZN(n18750) );
  INV_X1 U79 ( .A(n18770), .ZN(n18761) );
  INV_X1 U80 ( .A(n18781), .ZN(n18772) );
  INV_X1 U81 ( .A(n18792), .ZN(n18783) );
  INV_X1 U82 ( .A(n18803), .ZN(n18794) );
  INV_X1 U83 ( .A(n18814), .ZN(n18805) );
  INV_X1 U84 ( .A(n18825), .ZN(n18816) );
  INV_X1 U85 ( .A(n18836), .ZN(n18827) );
  INV_X1 U86 ( .A(n18847), .ZN(n18838) );
  INV_X1 U87 ( .A(n18858), .ZN(n18849) );
  INV_X1 U88 ( .A(n18869), .ZN(n18860) );
  INV_X1 U89 ( .A(n18880), .ZN(n18871) );
  INV_X1 U90 ( .A(n18891), .ZN(n18882) );
  INV_X1 U91 ( .A(n18902), .ZN(n18893) );
  INV_X1 U92 ( .A(n18989), .ZN(n18982) );
  INV_X1 U93 ( .A(n18571), .ZN(n18561) );
  INV_X1 U94 ( .A(n18585), .ZN(n18575) );
  INV_X1 U95 ( .A(n18611), .ZN(n18601) );
  INV_X1 U96 ( .A(n18658), .ZN(n18648) );
  INV_X1 U97 ( .A(n18749), .ZN(n18739) );
  INV_X1 U98 ( .A(n18571), .ZN(n18562) );
  INV_X1 U99 ( .A(n18585), .ZN(n18576) );
  INV_X1 U100 ( .A(n18611), .ZN(n18602) );
  INV_X1 U101 ( .A(n18658), .ZN(n18649) );
  INV_X1 U102 ( .A(n18749), .ZN(n18740) );
  BUF_X1 U103 ( .A(n18735), .Z(n18726) );
  BUF_X1 U104 ( .A(n18726), .Z(n18733) );
  BUF_X1 U105 ( .A(n18730), .Z(n18732) );
  BUF_X1 U106 ( .A(n18735), .Z(n18731) );
  BUF_X1 U107 ( .A(n18735), .Z(n18729) );
  BUF_X1 U108 ( .A(n18735), .Z(n18728) );
  BUF_X1 U109 ( .A(n18735), .Z(n18727) );
  BUF_X1 U110 ( .A(n18735), .Z(n18730) );
  BUF_X1 U111 ( .A(n18735), .Z(n18734) );
  NAND2_X1 U112 ( .A1(n4543), .A2(n4542), .ZN(n3949) );
  NAND2_X1 U113 ( .A1(n4543), .A2(n4539), .ZN(n3975) );
  NAND2_X1 U114 ( .A1(n4543), .A2(n4540), .ZN(n3980) );
  NAND2_X1 U115 ( .A1(n4532), .A2(n4539), .ZN(n3945) );
  NAND2_X1 U116 ( .A1(n4532), .A2(n4542), .ZN(n3969) );
  BUF_X1 U117 ( .A(n2213), .Z(n18502) );
  BUF_X1 U118 ( .A(n2213), .Z(n18503) );
  BUF_X1 U119 ( .A(n2218), .Z(n18499) );
  BUF_X1 U120 ( .A(n2218), .Z(n18500) );
  BUF_X1 U121 ( .A(n3965), .Z(n18395) );
  BUF_X1 U122 ( .A(n3965), .Z(n18396) );
  BUF_X1 U123 ( .A(n2220), .Z(n18493) );
  BUF_X1 U124 ( .A(n2222), .Z(n18487) );
  BUF_X1 U125 ( .A(n2235), .Z(n18454) );
  BUF_X1 U126 ( .A(n2230), .Z(n18466) );
  BUF_X1 U127 ( .A(n2220), .Z(n18494) );
  BUF_X1 U128 ( .A(n2222), .Z(n18488) );
  BUF_X1 U129 ( .A(n2235), .Z(n18455) );
  BUF_X1 U130 ( .A(n2230), .Z(n18467) );
  BUF_X1 U131 ( .A(n2219), .Z(n18496) );
  BUF_X1 U132 ( .A(n2236), .Z(n18451) );
  BUF_X1 U133 ( .A(n2219), .Z(n18497) );
  BUF_X1 U134 ( .A(n2236), .Z(n18452) );
  BUF_X1 U135 ( .A(n2231), .Z(n18463) );
  BUF_X1 U136 ( .A(n2231), .Z(n18464) );
  BUF_X1 U137 ( .A(n3968), .Z(n18386) );
  BUF_X1 U138 ( .A(n3966), .Z(n18392) );
  BUF_X1 U139 ( .A(n3968), .Z(n18387) );
  BUF_X1 U140 ( .A(n3966), .Z(n18393) );
  BUF_X1 U141 ( .A(n2221), .Z(n18490) );
  BUF_X1 U142 ( .A(n2223), .Z(n18484) );
  BUF_X1 U143 ( .A(n2221), .Z(n18491) );
  BUF_X1 U144 ( .A(n2223), .Z(n18485) );
  BUF_X1 U145 ( .A(n2205), .Z(n18520) );
  BUF_X1 U146 ( .A(n2205), .Z(n18521) );
  BUF_X1 U147 ( .A(n3955), .Z(n18410) );
  BUF_X1 U148 ( .A(n3950), .Z(n18422) );
  BUF_X1 U149 ( .A(n3955), .Z(n18411) );
  BUF_X1 U150 ( .A(n3950), .Z(n18423) );
  BUF_X1 U151 ( .A(n2200), .Z(n18532) );
  BUF_X1 U152 ( .A(n2195), .Z(n18543) );
  BUF_X1 U153 ( .A(n2210), .Z(n18508) );
  BUF_X1 U154 ( .A(n2200), .Z(n18533) );
  BUF_X1 U155 ( .A(n2195), .Z(n18544) );
  BUF_X1 U156 ( .A(n2210), .Z(n18509) );
  BUF_X1 U157 ( .A(n2232), .Z(n18460) );
  BUF_X1 U158 ( .A(n2227), .Z(n18472) );
  BUF_X1 U159 ( .A(n2232), .Z(n18461) );
  BUF_X1 U160 ( .A(n2227), .Z(n18473) );
  BUF_X1 U161 ( .A(n3972), .Z(n18374) );
  BUF_X1 U162 ( .A(n3972), .Z(n18375) );
  BUF_X1 U163 ( .A(n2197), .Z(n18540) );
  BUF_X1 U164 ( .A(n2197), .Z(n18541) );
  BUF_X1 U165 ( .A(n3952), .Z(n18419) );
  BUF_X1 U166 ( .A(n3947), .Z(n18431) );
  BUF_X1 U167 ( .A(n3952), .Z(n18420) );
  BUF_X1 U168 ( .A(n3947), .Z(n18432) );
  BUF_X1 U169 ( .A(n2202), .Z(n18529) );
  BUF_X1 U170 ( .A(n2207), .Z(n18517) );
  BUF_X1 U171 ( .A(n2212), .Z(n18505) );
  BUF_X1 U172 ( .A(n2202), .Z(n18530) );
  BUF_X1 U173 ( .A(n2207), .Z(n18518) );
  BUF_X1 U174 ( .A(n2212), .Z(n18506) );
  BUF_X1 U175 ( .A(n2233), .Z(n18457) );
  BUF_X1 U176 ( .A(n2233), .Z(n18458) );
  BUF_X1 U177 ( .A(n3973), .Z(n18371) );
  BUF_X1 U178 ( .A(n3973), .Z(n18372) );
  BUF_X1 U179 ( .A(n2228), .Z(n18469) );
  BUF_X1 U180 ( .A(n2228), .Z(n18470) );
  BUF_X1 U181 ( .A(n2204), .Z(n18523) );
  BUF_X1 U182 ( .A(n2204), .Z(n18524) );
  BUF_X1 U183 ( .A(n2199), .Z(n18535) );
  BUF_X1 U184 ( .A(n2194), .Z(n18546) );
  BUF_X1 U185 ( .A(n2209), .Z(n18511) );
  BUF_X1 U186 ( .A(n2199), .Z(n18536) );
  BUF_X1 U187 ( .A(n2194), .Z(n18547) );
  BUF_X1 U188 ( .A(n2209), .Z(n18512) );
  BUF_X1 U189 ( .A(n3954), .Z(n18413) );
  BUF_X1 U190 ( .A(n3939), .Z(n18448) );
  BUF_X1 U191 ( .A(n3944), .Z(n18437) );
  BUF_X1 U192 ( .A(n3954), .Z(n18414) );
  BUF_X1 U193 ( .A(n3939), .Z(n18449) );
  BUF_X1 U194 ( .A(n3944), .Z(n18438) );
  BUF_X1 U195 ( .A(n2226), .Z(n18475) );
  BUF_X1 U196 ( .A(n2226), .Z(n18476) );
  BUF_X1 U197 ( .A(n3971), .Z(n18377) );
  BUF_X1 U198 ( .A(n3971), .Z(n18378) );
  BUF_X1 U199 ( .A(n2218), .Z(n18501) );
  BUF_X1 U200 ( .A(n3965), .Z(n18397) );
  BUF_X1 U201 ( .A(n2220), .Z(n18495) );
  BUF_X1 U202 ( .A(n2222), .Z(n18489) );
  BUF_X1 U203 ( .A(n2235), .Z(n18456) );
  BUF_X1 U204 ( .A(n2230), .Z(n18468) );
  BUF_X1 U205 ( .A(n2213), .Z(n18504) );
  BUF_X1 U206 ( .A(n2224), .Z(n18481) );
  BUF_X1 U207 ( .A(n2224), .Z(n18482) );
  BUF_X1 U208 ( .A(n3970), .Z(n18380) );
  BUF_X1 U209 ( .A(n3970), .Z(n18381) );
  BUF_X1 U210 ( .A(n2225), .Z(n18478) );
  BUF_X1 U211 ( .A(n2225), .Z(n18479) );
  BUF_X1 U212 ( .A(n2219), .Z(n18498) );
  BUF_X1 U213 ( .A(n2236), .Z(n18453) );
  BUF_X1 U214 ( .A(n2231), .Z(n18465) );
  BUF_X1 U215 ( .A(n3968), .Z(n18388) );
  BUF_X1 U216 ( .A(n3966), .Z(n18394) );
  BUF_X1 U217 ( .A(n2221), .Z(n18492) );
  BUF_X1 U218 ( .A(n2223), .Z(n18486) );
  BUF_X1 U219 ( .A(n2203), .Z(n18527) );
  BUF_X1 U220 ( .A(n2208), .Z(n18515) );
  BUF_X1 U221 ( .A(n2203), .Z(n18526) );
  BUF_X1 U222 ( .A(n2208), .Z(n18514) );
  BUF_X1 U223 ( .A(n3953), .Z(n18417) );
  BUF_X1 U224 ( .A(n3948), .Z(n18429) );
  BUF_X1 U225 ( .A(n3953), .Z(n18416) );
  BUF_X1 U226 ( .A(n3948), .Z(n18428) );
  BUF_X1 U227 ( .A(n2205), .Z(n18522) );
  BUF_X1 U228 ( .A(n3955), .Z(n18412) );
  BUF_X1 U229 ( .A(n3950), .Z(n18424) );
  BUF_X1 U230 ( .A(n2200), .Z(n18534) );
  BUF_X1 U231 ( .A(n2195), .Z(n18545) );
  BUF_X1 U232 ( .A(n2210), .Z(n18510) );
  BUF_X1 U233 ( .A(n2232), .Z(n18462) );
  BUF_X1 U234 ( .A(n2227), .Z(n18474) );
  BUF_X1 U235 ( .A(n3972), .Z(n18376) );
  BUF_X1 U236 ( .A(n2197), .Z(n18542) );
  BUF_X1 U237 ( .A(n3952), .Z(n18421) );
  BUF_X1 U238 ( .A(n3947), .Z(n18433) );
  BUF_X1 U239 ( .A(n2202), .Z(n18531) );
  BUF_X1 U240 ( .A(n2207), .Z(n18519) );
  BUF_X1 U241 ( .A(n2212), .Z(n18507) );
  BUF_X1 U242 ( .A(n2233), .Z(n18459) );
  BUF_X1 U243 ( .A(n3973), .Z(n18373) );
  BUF_X1 U244 ( .A(n2228), .Z(n18471) );
  BUF_X1 U245 ( .A(n2204), .Z(n18525) );
  BUF_X1 U246 ( .A(n2199), .Z(n18537) );
  BUF_X1 U247 ( .A(n2194), .Z(n18548) );
  BUF_X1 U248 ( .A(n2209), .Z(n18513) );
  BUF_X1 U249 ( .A(n3954), .Z(n18415) );
  BUF_X1 U250 ( .A(n3939), .Z(n18450) );
  BUF_X1 U251 ( .A(n3944), .Z(n18439) );
  BUF_X1 U252 ( .A(n2226), .Z(n18477) );
  BUF_X1 U253 ( .A(n3971), .Z(n18379) );
  BUF_X1 U254 ( .A(n2224), .Z(n18483) );
  BUF_X1 U255 ( .A(n3970), .Z(n18382) );
  BUF_X1 U256 ( .A(n2225), .Z(n18480) );
  BUF_X1 U257 ( .A(n2203), .Z(n18528) );
  BUF_X1 U258 ( .A(n2208), .Z(n18516) );
  BUF_X1 U259 ( .A(n3953), .Z(n18418) );
  BUF_X1 U260 ( .A(n3948), .Z(n18430) );
  NAND2_X1 U261 ( .A1(n4537), .A2(n4543), .ZN(n3976) );
  NAND2_X1 U262 ( .A1(n4545), .A2(n4543), .ZN(n3963) );
  NAND2_X1 U263 ( .A1(n4533), .A2(n4543), .ZN(n3967) );
  NAND2_X1 U264 ( .A1(n4533), .A2(n4532), .ZN(n3940) );
  NAND2_X1 U265 ( .A1(n4545), .A2(n4532), .ZN(n3964) );
  NAND2_X1 U266 ( .A1(n4534), .A2(n4532), .ZN(n3981) );
  AND2_X1 U267 ( .A1(n4543), .A2(n4531), .ZN(n3978) );
  AND2_X1 U268 ( .A1(n4534), .A2(n4543), .ZN(n3957) );
  AND2_X1 U269 ( .A1(n4540), .A2(n4532), .ZN(n3958) );
  AND2_X1 U270 ( .A1(n4531), .A2(n4532), .ZN(n3942) );
  AND2_X1 U271 ( .A1(n4537), .A2(n4532), .ZN(n3977) );
  INV_X1 U272 ( .A(n18557), .ZN(n18550) );
  INV_X1 U273 ( .A(n18557), .ZN(n18549) );
  BUF_X1 U274 ( .A(n18990), .Z(n18983) );
  BUF_X1 U275 ( .A(n18990), .Z(n18984) );
  BUF_X1 U276 ( .A(n18990), .Z(n18985) );
  BUF_X1 U277 ( .A(n18990), .Z(n18986) );
  BUF_X1 U278 ( .A(n18990), .Z(n18987) );
  BUF_X1 U279 ( .A(n18990), .Z(n18988) );
  BUF_X1 U280 ( .A(n18990), .Z(n18989) );
  BUF_X1 U281 ( .A(n18560), .Z(n18571) );
  BUF_X1 U282 ( .A(n18574), .Z(n18585) );
  BUF_X1 U283 ( .A(n18600), .Z(n18611) );
  BUF_X1 U284 ( .A(n18647), .Z(n18658) );
  BUF_X1 U285 ( .A(n18738), .Z(n18749) );
  BUF_X1 U286 ( .A(n18597), .Z(n18588) );
  BUF_X1 U287 ( .A(n18622), .Z(n18613) );
  BUF_X1 U288 ( .A(n18633), .Z(n18624) );
  BUF_X1 U289 ( .A(n18669), .Z(n18660) );
  BUF_X1 U290 ( .A(n18680), .Z(n18671) );
  BUF_X1 U291 ( .A(n18702), .Z(n18693) );
  BUF_X1 U292 ( .A(n18760), .Z(n18751) );
  BUF_X1 U293 ( .A(n18771), .Z(n18762) );
  BUF_X1 U294 ( .A(n18793), .Z(n18784) );
  BUF_X1 U295 ( .A(n18837), .Z(n18828) );
  BUF_X1 U296 ( .A(n18644), .Z(n18635) );
  BUF_X1 U297 ( .A(n18691), .Z(n18682) );
  BUF_X1 U298 ( .A(n18713), .Z(n18704) );
  BUF_X1 U299 ( .A(n18724), .Z(n18715) );
  BUF_X1 U300 ( .A(n18782), .Z(n18773) );
  BUF_X1 U301 ( .A(n18804), .Z(n18795) );
  BUF_X1 U302 ( .A(n18815), .Z(n18806) );
  BUF_X1 U303 ( .A(n18848), .Z(n18839) );
  BUF_X1 U304 ( .A(n18859), .Z(n18850) );
  BUF_X1 U305 ( .A(n18881), .Z(n18872) );
  BUF_X1 U306 ( .A(n18826), .Z(n18817) );
  BUF_X1 U307 ( .A(n18870), .Z(n18861) );
  BUF_X1 U308 ( .A(n18892), .Z(n18883) );
  BUF_X1 U309 ( .A(n18903), .Z(n18894) );
  BUF_X1 U310 ( .A(n18560), .Z(n18569) );
  BUF_X1 U311 ( .A(n18559), .Z(n18568) );
  BUF_X1 U312 ( .A(n18559), .Z(n18567) );
  BUF_X1 U313 ( .A(n18559), .Z(n18566) );
  BUF_X1 U314 ( .A(n18558), .Z(n18565) );
  BUF_X1 U315 ( .A(n18558), .Z(n18564) );
  BUF_X1 U316 ( .A(n18558), .Z(n18563) );
  BUF_X1 U317 ( .A(n18574), .Z(n18583) );
  BUF_X1 U318 ( .A(n18573), .Z(n18582) );
  BUF_X1 U319 ( .A(n18573), .Z(n18580) );
  BUF_X1 U320 ( .A(n18572), .Z(n18579) );
  BUF_X1 U321 ( .A(n18572), .Z(n18578) );
  BUF_X1 U322 ( .A(n18572), .Z(n18577) );
  BUF_X1 U323 ( .A(n18573), .Z(n18581) );
  BUF_X1 U324 ( .A(n18600), .Z(n18609) );
  BUF_X1 U325 ( .A(n18599), .Z(n18608) );
  BUF_X1 U326 ( .A(n18599), .Z(n18606) );
  BUF_X1 U327 ( .A(n18598), .Z(n18605) );
  BUF_X1 U328 ( .A(n18598), .Z(n18604) );
  BUF_X1 U329 ( .A(n18598), .Z(n18603) );
  BUF_X1 U330 ( .A(n18599), .Z(n18607) );
  BUF_X1 U331 ( .A(n18647), .Z(n18656) );
  BUF_X1 U332 ( .A(n18646), .Z(n18655) );
  BUF_X1 U333 ( .A(n18646), .Z(n18653) );
  BUF_X1 U334 ( .A(n18645), .Z(n18652) );
  BUF_X1 U335 ( .A(n18645), .Z(n18651) );
  BUF_X1 U336 ( .A(n18645), .Z(n18650) );
  BUF_X1 U337 ( .A(n18646), .Z(n18654) );
  BUF_X1 U338 ( .A(n18738), .Z(n18747) );
  BUF_X1 U339 ( .A(n18737), .Z(n18746) );
  BUF_X1 U340 ( .A(n18737), .Z(n18744) );
  BUF_X1 U341 ( .A(n18736), .Z(n18743) );
  BUF_X1 U342 ( .A(n18736), .Z(n18742) );
  BUF_X1 U343 ( .A(n18736), .Z(n18741) );
  BUF_X1 U344 ( .A(n18737), .Z(n18745) );
  BUF_X1 U345 ( .A(n18560), .Z(n18570) );
  BUF_X1 U346 ( .A(n18574), .Z(n18584) );
  BUF_X1 U347 ( .A(n18600), .Z(n18610) );
  BUF_X1 U348 ( .A(n18647), .Z(n18657) );
  BUF_X1 U349 ( .A(n18738), .Z(n18748) );
  BUF_X1 U350 ( .A(n18588), .Z(n18595) );
  BUF_X1 U351 ( .A(n18592), .Z(n18594) );
  BUF_X1 U352 ( .A(n18597), .Z(n18593) );
  BUF_X1 U353 ( .A(n18597), .Z(n18591) );
  BUF_X1 U354 ( .A(n18597), .Z(n18590) );
  BUF_X1 U355 ( .A(n18597), .Z(n18589) );
  BUF_X1 U356 ( .A(n18597), .Z(n18592) );
  BUF_X1 U357 ( .A(n18613), .Z(n18620) );
  BUF_X1 U358 ( .A(n18617), .Z(n18619) );
  BUF_X1 U359 ( .A(n18622), .Z(n18618) );
  BUF_X1 U360 ( .A(n18622), .Z(n18616) );
  BUF_X1 U361 ( .A(n18622), .Z(n18615) );
  BUF_X1 U362 ( .A(n18622), .Z(n18614) );
  BUF_X1 U363 ( .A(n18622), .Z(n18617) );
  BUF_X1 U364 ( .A(n18624), .Z(n18631) );
  BUF_X1 U365 ( .A(n18625), .Z(n18630) );
  BUF_X1 U366 ( .A(n18633), .Z(n18629) );
  BUF_X1 U367 ( .A(n18633), .Z(n18627) );
  BUF_X1 U368 ( .A(n18633), .Z(n18626) );
  BUF_X1 U369 ( .A(n18633), .Z(n18625) );
  BUF_X1 U370 ( .A(n18633), .Z(n18628) );
  BUF_X1 U371 ( .A(n18635), .Z(n18642) );
  BUF_X1 U372 ( .A(n18639), .Z(n18641) );
  BUF_X1 U373 ( .A(n18644), .Z(n18640) );
  BUF_X1 U374 ( .A(n18644), .Z(n18638) );
  BUF_X1 U375 ( .A(n18644), .Z(n18637) );
  BUF_X1 U376 ( .A(n18644), .Z(n18636) );
  BUF_X1 U377 ( .A(n18644), .Z(n18639) );
  BUF_X1 U378 ( .A(n18660), .Z(n18667) );
  BUF_X1 U379 ( .A(n18664), .Z(n18666) );
  BUF_X1 U380 ( .A(n18669), .Z(n18665) );
  BUF_X1 U381 ( .A(n18669), .Z(n18663) );
  BUF_X1 U382 ( .A(n18669), .Z(n18662) );
  BUF_X1 U383 ( .A(n18669), .Z(n18661) );
  BUF_X1 U384 ( .A(n18669), .Z(n18664) );
  BUF_X1 U385 ( .A(n18671), .Z(n18678) );
  BUF_X1 U386 ( .A(n18675), .Z(n18677) );
  BUF_X1 U387 ( .A(n18680), .Z(n18676) );
  BUF_X1 U388 ( .A(n18680), .Z(n18674) );
  BUF_X1 U389 ( .A(n18680), .Z(n18673) );
  BUF_X1 U390 ( .A(n18680), .Z(n18672) );
  BUF_X1 U391 ( .A(n18680), .Z(n18675) );
  BUF_X1 U392 ( .A(n18682), .Z(n18689) );
  BUF_X1 U393 ( .A(n18686), .Z(n18688) );
  BUF_X1 U394 ( .A(n18691), .Z(n18687) );
  BUF_X1 U395 ( .A(n18691), .Z(n18685) );
  BUF_X1 U396 ( .A(n18691), .Z(n18684) );
  BUF_X1 U397 ( .A(n18691), .Z(n18683) );
  BUF_X1 U398 ( .A(n18691), .Z(n18686) );
  BUF_X1 U399 ( .A(n18693), .Z(n18700) );
  BUF_X1 U400 ( .A(n18697), .Z(n18699) );
  BUF_X1 U401 ( .A(n18702), .Z(n18698) );
  BUF_X1 U402 ( .A(n18702), .Z(n18696) );
  BUF_X1 U403 ( .A(n18702), .Z(n18695) );
  BUF_X1 U404 ( .A(n18702), .Z(n18694) );
  BUF_X1 U405 ( .A(n18702), .Z(n18697) );
  BUF_X1 U406 ( .A(n18704), .Z(n18711) );
  BUF_X1 U407 ( .A(n18708), .Z(n18710) );
  BUF_X1 U408 ( .A(n18713), .Z(n18709) );
  BUF_X1 U409 ( .A(n18713), .Z(n18707) );
  BUF_X1 U410 ( .A(n18713), .Z(n18706) );
  BUF_X1 U411 ( .A(n18713), .Z(n18705) );
  BUF_X1 U412 ( .A(n18713), .Z(n18708) );
  BUF_X1 U413 ( .A(n18715), .Z(n18722) );
  BUF_X1 U414 ( .A(n18719), .Z(n18721) );
  BUF_X1 U415 ( .A(n18724), .Z(n18720) );
  BUF_X1 U416 ( .A(n18724), .Z(n18718) );
  BUF_X1 U417 ( .A(n18724), .Z(n18717) );
  BUF_X1 U418 ( .A(n18724), .Z(n18716) );
  BUF_X1 U419 ( .A(n18724), .Z(n18719) );
  BUF_X1 U420 ( .A(n18751), .Z(n18758) );
  BUF_X1 U421 ( .A(n18755), .Z(n18757) );
  BUF_X1 U422 ( .A(n18760), .Z(n18756) );
  BUF_X1 U423 ( .A(n18760), .Z(n18754) );
  BUF_X1 U424 ( .A(n18760), .Z(n18753) );
  BUF_X1 U425 ( .A(n18760), .Z(n18752) );
  BUF_X1 U426 ( .A(n18760), .Z(n18755) );
  BUF_X1 U427 ( .A(n18762), .Z(n18769) );
  BUF_X1 U428 ( .A(n18766), .Z(n18768) );
  BUF_X1 U429 ( .A(n18771), .Z(n18767) );
  BUF_X1 U430 ( .A(n18771), .Z(n18765) );
  BUF_X1 U431 ( .A(n18771), .Z(n18764) );
  BUF_X1 U432 ( .A(n18771), .Z(n18763) );
  BUF_X1 U433 ( .A(n18771), .Z(n18766) );
  BUF_X1 U434 ( .A(n18773), .Z(n18780) );
  BUF_X1 U435 ( .A(n18777), .Z(n18779) );
  BUF_X1 U436 ( .A(n18782), .Z(n18778) );
  BUF_X1 U437 ( .A(n18782), .Z(n18776) );
  BUF_X1 U438 ( .A(n18782), .Z(n18775) );
  BUF_X1 U439 ( .A(n18782), .Z(n18774) );
  BUF_X1 U440 ( .A(n18782), .Z(n18777) );
  BUF_X1 U441 ( .A(n18784), .Z(n18791) );
  BUF_X1 U442 ( .A(n18788), .Z(n18790) );
  BUF_X1 U443 ( .A(n18793), .Z(n18789) );
  BUF_X1 U444 ( .A(n18793), .Z(n18787) );
  BUF_X1 U445 ( .A(n18793), .Z(n18786) );
  BUF_X1 U446 ( .A(n18793), .Z(n18785) );
  BUF_X1 U447 ( .A(n18793), .Z(n18788) );
  BUF_X1 U448 ( .A(n18795), .Z(n18802) );
  BUF_X1 U449 ( .A(n18799), .Z(n18801) );
  BUF_X1 U450 ( .A(n18804), .Z(n18800) );
  BUF_X1 U451 ( .A(n18804), .Z(n18798) );
  BUF_X1 U452 ( .A(n18804), .Z(n18797) );
  BUF_X1 U453 ( .A(n18804), .Z(n18796) );
  BUF_X1 U454 ( .A(n18804), .Z(n18799) );
  BUF_X1 U455 ( .A(n18806), .Z(n18813) );
  BUF_X1 U456 ( .A(n18810), .Z(n18812) );
  BUF_X1 U457 ( .A(n18815), .Z(n18811) );
  BUF_X1 U458 ( .A(n18815), .Z(n18809) );
  BUF_X1 U459 ( .A(n18815), .Z(n18808) );
  BUF_X1 U460 ( .A(n18815), .Z(n18807) );
  BUF_X1 U461 ( .A(n18815), .Z(n18810) );
  BUF_X1 U462 ( .A(n18817), .Z(n18824) );
  BUF_X1 U463 ( .A(n18821), .Z(n18823) );
  BUF_X1 U464 ( .A(n18826), .Z(n18822) );
  BUF_X1 U465 ( .A(n18826), .Z(n18820) );
  BUF_X1 U466 ( .A(n18826), .Z(n18819) );
  BUF_X1 U467 ( .A(n18826), .Z(n18818) );
  BUF_X1 U468 ( .A(n18826), .Z(n18821) );
  BUF_X1 U469 ( .A(n18837), .Z(n18829) );
  BUF_X1 U470 ( .A(n18837), .Z(n18830) );
  BUF_X1 U471 ( .A(n18837), .Z(n18831) );
  BUF_X1 U472 ( .A(n18837), .Z(n18832) );
  BUF_X1 U473 ( .A(n18837), .Z(n18833) );
  BUF_X1 U474 ( .A(n18829), .Z(n18834) );
  BUF_X1 U475 ( .A(n18828), .Z(n18835) );
  BUF_X1 U476 ( .A(n18839), .Z(n18846) );
  BUF_X1 U477 ( .A(n18843), .Z(n18845) );
  BUF_X1 U478 ( .A(n18848), .Z(n18844) );
  BUF_X1 U479 ( .A(n18848), .Z(n18842) );
  BUF_X1 U480 ( .A(n18848), .Z(n18841) );
  BUF_X1 U481 ( .A(n18848), .Z(n18840) );
  BUF_X1 U482 ( .A(n18848), .Z(n18843) );
  BUF_X1 U483 ( .A(n18850), .Z(n18857) );
  BUF_X1 U484 ( .A(n18854), .Z(n18856) );
  BUF_X1 U485 ( .A(n18859), .Z(n18855) );
  BUF_X1 U486 ( .A(n18859), .Z(n18853) );
  BUF_X1 U487 ( .A(n18859), .Z(n18852) );
  BUF_X1 U488 ( .A(n18859), .Z(n18851) );
  BUF_X1 U489 ( .A(n18859), .Z(n18854) );
  BUF_X1 U490 ( .A(n18861), .Z(n18868) );
  BUF_X1 U491 ( .A(n18865), .Z(n18867) );
  BUF_X1 U492 ( .A(n18870), .Z(n18866) );
  BUF_X1 U493 ( .A(n18870), .Z(n18864) );
  BUF_X1 U494 ( .A(n18870), .Z(n18863) );
  BUF_X1 U495 ( .A(n18870), .Z(n18862) );
  BUF_X1 U496 ( .A(n18870), .Z(n18865) );
  BUF_X1 U497 ( .A(n18881), .Z(n18873) );
  BUF_X1 U498 ( .A(n18881), .Z(n18874) );
  BUF_X1 U499 ( .A(n18881), .Z(n18875) );
  BUF_X1 U500 ( .A(n18881), .Z(n18876) );
  BUF_X1 U501 ( .A(n18881), .Z(n18877) );
  BUF_X1 U502 ( .A(n18873), .Z(n18878) );
  BUF_X1 U503 ( .A(n18872), .Z(n18879) );
  BUF_X1 U504 ( .A(n18883), .Z(n18890) );
  BUF_X1 U505 ( .A(n18887), .Z(n18889) );
  BUF_X1 U506 ( .A(n18892), .Z(n18888) );
  BUF_X1 U507 ( .A(n18892), .Z(n18886) );
  BUF_X1 U508 ( .A(n18892), .Z(n18885) );
  BUF_X1 U509 ( .A(n18892), .Z(n18884) );
  BUF_X1 U510 ( .A(n18892), .Z(n18887) );
  BUF_X1 U511 ( .A(n18903), .Z(n18895) );
  BUF_X1 U512 ( .A(n18903), .Z(n18896) );
  BUF_X1 U513 ( .A(n18903), .Z(n18897) );
  BUF_X1 U514 ( .A(n18903), .Z(n18898) );
  BUF_X1 U515 ( .A(n18903), .Z(n18899) );
  BUF_X1 U516 ( .A(n18895), .Z(n18900) );
  BUF_X1 U517 ( .A(n18894), .Z(n18901) );
  BUF_X1 U518 ( .A(n18597), .Z(n18596) );
  BUF_X1 U519 ( .A(n18622), .Z(n18621) );
  BUF_X1 U520 ( .A(n18633), .Z(n18632) );
  BUF_X1 U521 ( .A(n18644), .Z(n18643) );
  BUF_X1 U522 ( .A(n18669), .Z(n18668) );
  BUF_X1 U523 ( .A(n18680), .Z(n18679) );
  BUF_X1 U524 ( .A(n18691), .Z(n18690) );
  BUF_X1 U525 ( .A(n18702), .Z(n18701) );
  BUF_X1 U526 ( .A(n18713), .Z(n18712) );
  BUF_X1 U527 ( .A(n18724), .Z(n18723) );
  BUF_X1 U528 ( .A(n18760), .Z(n18759) );
  BUF_X1 U529 ( .A(n18771), .Z(n18770) );
  BUF_X1 U530 ( .A(n18782), .Z(n18781) );
  BUF_X1 U531 ( .A(n18793), .Z(n18792) );
  BUF_X1 U532 ( .A(n18804), .Z(n18803) );
  BUF_X1 U533 ( .A(n18815), .Z(n18814) );
  BUF_X1 U534 ( .A(n18826), .Z(n18825) );
  BUF_X1 U535 ( .A(n18837), .Z(n18836) );
  BUF_X1 U536 ( .A(n18848), .Z(n18847) );
  BUF_X1 U537 ( .A(n18859), .Z(n18858) );
  BUF_X1 U538 ( .A(n18870), .Z(n18869) );
  BUF_X1 U539 ( .A(n18881), .Z(n18880) );
  BUF_X1 U540 ( .A(n18892), .Z(n18891) );
  BUF_X1 U541 ( .A(n18903), .Z(n18902) );
  INV_X1 U542 ( .A(n1666), .ZN(n18735) );
  NOR3_X1 U543 ( .A1(n3929), .A2(n3926), .A3(n3928), .ZN(n3919) );
  NAND2_X1 U544 ( .A1(n3917), .A2(n3912), .ZN(n2218) );
  NAND2_X1 U545 ( .A1(n3906), .A2(n3915), .ZN(n2199) );
  NAND2_X1 U546 ( .A1(n3906), .A2(n3909), .ZN(n2194) );
  NAND2_X1 U547 ( .A1(n3906), .A2(n3908), .ZN(n2209) );
  NAND2_X1 U548 ( .A1(n3906), .A2(n3913), .ZN(n2231) );
  NAND2_X1 U549 ( .A1(n3909), .A2(n3917), .ZN(n2204) );
  NAND2_X1 U550 ( .A1(n3905), .A2(n3917), .ZN(n2205) );
  NAND2_X1 U551 ( .A1(n3911), .A2(n3917), .ZN(n2226) );
  NAND2_X1 U552 ( .A1(n3919), .A2(n3917), .ZN(n2219) );
  NAND2_X1 U553 ( .A1(n3913), .A2(n3917), .ZN(n2236) );
  NAND2_X1 U554 ( .A1(n3909), .A2(n3907), .ZN(n2222) );
  NAND2_X1 U555 ( .A1(n3909), .A2(n3914), .ZN(n2235) );
  NAND2_X1 U556 ( .A1(n3908), .A2(n3914), .ZN(n2224) );
  NAND2_X1 U557 ( .A1(n3911), .A2(n3914), .ZN(n2221) );
  NAND2_X1 U558 ( .A1(n4540), .A2(n4535), .ZN(n3944) );
  NAND2_X1 U559 ( .A1(n4540), .A2(n4538), .ZN(n3968) );
  NAND2_X1 U560 ( .A1(n3913), .A2(n3914), .ZN(n2200) );
  NAND2_X1 U561 ( .A1(n3912), .A2(n3914), .ZN(n2225) );
  NAND2_X1 U562 ( .A1(n4531), .A2(n4538), .ZN(n3971) );
  NAND2_X1 U563 ( .A1(n4531), .A2(n4535), .ZN(n3966) );
  NAND2_X1 U564 ( .A1(n3919), .A2(n3907), .ZN(n2220) );
  NAND2_X1 U565 ( .A1(n4534), .A2(n4535), .ZN(n3939) );
  NAND2_X1 U566 ( .A1(n3905), .A2(n3914), .ZN(n2230) );
  NAND2_X1 U567 ( .A1(n3907), .A2(n3908), .ZN(n2195) );
  NAND2_X1 U568 ( .A1(n3907), .A2(n3911), .ZN(n2210) );
  NAND2_X1 U569 ( .A1(n3907), .A2(n3915), .ZN(n2223) );
  AND2_X1 U570 ( .A1(n3917), .A2(n3908), .ZN(n2227) );
  NAND2_X1 U571 ( .A1(n4535), .A2(n4539), .ZN(n3970) );
  AND2_X1 U572 ( .A1(n3906), .A2(n3911), .ZN(n2203) );
  AND2_X1 U573 ( .A1(n3906), .A2(n3912), .ZN(n2208) );
  AND2_X1 U574 ( .A1(n3906), .A2(n3919), .ZN(n2232) );
  NAND2_X1 U575 ( .A1(n4533), .A2(n4535), .ZN(n3950) );
  NAND2_X1 U576 ( .A1(n4545), .A2(n4535), .ZN(n3965) );
  AND2_X1 U577 ( .A1(n3915), .A2(n3917), .ZN(n2233) );
  NAND2_X1 U578 ( .A1(n4545), .A2(n4538), .ZN(n3955) );
  NAND2_X1 U579 ( .A1(n4538), .A2(n4539), .ZN(n3954) );
  AND2_X1 U580 ( .A1(n3905), .A2(n3906), .ZN(n2197) );
  AND2_X1 U581 ( .A1(n3913), .A2(n3907), .ZN(n2212) );
  AND2_X1 U582 ( .A1(n3915), .A2(n3914), .ZN(n2228) );
  AND2_X1 U583 ( .A1(n3919), .A2(n3914), .ZN(n2213) );
  AND2_X1 U584 ( .A1(n4534), .A2(n4538), .ZN(n3947) );
  AND2_X1 U585 ( .A1(n3905), .A2(n3907), .ZN(n2207) );
  AND2_X1 U586 ( .A1(n4537), .A2(n4535), .ZN(n3952) );
  AND2_X1 U587 ( .A1(n4537), .A2(n4538), .ZN(n3948) );
  AND2_X1 U588 ( .A1(n3907), .A2(n3912), .ZN(n2202) );
  AND2_X1 U589 ( .A1(n4538), .A2(n4542), .ZN(n3972) );
  AND2_X1 U590 ( .A1(n4542), .A2(n4535), .ZN(n3953) );
  AND2_X1 U591 ( .A1(n4533), .A2(n4538), .ZN(n3973) );
  NOR3_X1 U592 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(ADD_RD2[0]), .ZN(n4540)
         );
  INV_X1 U593 ( .A(n18996), .ZN(n18999) );
  INV_X1 U594 ( .A(n18996), .ZN(n18998) );
  INV_X1 U595 ( .A(n18996), .ZN(n18997) );
  NOR3_X1 U596 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(n4550), .ZN(n4531) );
  NOR3_X1 U597 ( .A1(n4551), .A2(ADD_RD2[3]), .A3(n4550), .ZN(n4534) );
  NOR3_X1 U598 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[3]), .A3(n4551), .ZN(n4537) );
  AND3_X1 U599 ( .A1(ADD_RD2[3]), .A2(n4550), .A3(ADD_RD2[4]), .ZN(n4539) );
  AND3_X1 U600 ( .A1(n4550), .A2(n4551), .A3(ADD_RD2[3]), .ZN(n4545) );
  AND3_X1 U601 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .A3(ADD_RD2[0]), .ZN(n4533)
         );
  AND3_X1 U602 ( .A1(ADD_RD2[3]), .A2(n4551), .A3(ADD_RD2[0]), .ZN(n4542) );
  BUF_X1 U603 ( .A(n2183), .Z(n18556) );
  BUF_X1 U604 ( .A(n2183), .Z(n18555) );
  BUF_X1 U605 ( .A(n2183), .Z(n18554) );
  BUF_X1 U606 ( .A(n2183), .Z(n18553) );
  BUF_X1 U607 ( .A(n2183), .Z(n18552) );
  BUF_X1 U608 ( .A(n2183), .Z(n18551) );
  BUF_X1 U609 ( .A(n2183), .Z(n18557) );
  INV_X1 U610 ( .A(ADD_RD2[0]), .ZN(n4550) );
  INV_X1 U611 ( .A(ADD_RD2[4]), .ZN(n4551) );
  OAI21_X1 U612 ( .B1(n1139), .B2(n1700), .A(n18999), .ZN(n1666) );
  INV_X1 U613 ( .A(n1074), .ZN(n18990) );
  OAI21_X1 U614 ( .B1(n1138), .B2(n1139), .A(n18998), .ZN(n1074) );
  INV_X1 U615 ( .A(ADD_RD2[2]), .ZN(n4553) );
  BUF_X1 U616 ( .A(n2150), .Z(n18560) );
  BUF_X1 U617 ( .A(n2116), .Z(n18574) );
  BUF_X1 U618 ( .A(n2045), .Z(n18600) );
  BUF_X1 U619 ( .A(n1908), .Z(n18647) );
  BUF_X1 U620 ( .A(n1631), .Z(n18738) );
  BUF_X1 U621 ( .A(n2150), .Z(n18559) );
  BUF_X1 U622 ( .A(n2150), .Z(n18558) );
  BUF_X1 U623 ( .A(n2116), .Z(n18572) );
  BUF_X1 U624 ( .A(n2116), .Z(n18573) );
  BUF_X1 U625 ( .A(n2045), .Z(n18598) );
  BUF_X1 U626 ( .A(n2045), .Z(n18599) );
  BUF_X1 U627 ( .A(n1908), .Z(n18645) );
  BUF_X1 U628 ( .A(n1908), .Z(n18646) );
  BUF_X1 U629 ( .A(n1631), .Z(n18736) );
  BUF_X1 U630 ( .A(n1631), .Z(n18737) );
  INV_X1 U631 ( .A(n2079), .ZN(n18597) );
  INV_X1 U632 ( .A(n2011), .ZN(n18622) );
  INV_X1 U633 ( .A(n1977), .ZN(n18633) );
  INV_X1 U634 ( .A(n1942), .ZN(n18644) );
  INV_X1 U635 ( .A(n1874), .ZN(n18669) );
  INV_X1 U636 ( .A(n1840), .ZN(n18680) );
  INV_X1 U637 ( .A(n1805), .ZN(n18691) );
  INV_X1 U638 ( .A(n1770), .ZN(n18702) );
  INV_X1 U639 ( .A(n1736), .ZN(n18713) );
  INV_X1 U640 ( .A(n1702), .ZN(n18724) );
  INV_X1 U641 ( .A(n1597), .ZN(n18760) );
  INV_X1 U642 ( .A(n1563), .ZN(n18771) );
  INV_X1 U643 ( .A(n1528), .ZN(n18782) );
  INV_X1 U644 ( .A(n1494), .ZN(n18793) );
  INV_X1 U645 ( .A(n1460), .ZN(n18804) );
  INV_X1 U646 ( .A(n1426), .ZN(n18815) );
  INV_X1 U647 ( .A(n1390), .ZN(n18826) );
  INV_X1 U648 ( .A(n1356), .ZN(n18837) );
  INV_X1 U649 ( .A(n1322), .ZN(n18848) );
  INV_X1 U650 ( .A(n1288), .ZN(n18859) );
  INV_X1 U651 ( .A(n1252), .ZN(n18870) );
  INV_X1 U652 ( .A(n1214), .ZN(n18881) );
  INV_X1 U653 ( .A(n1178), .ZN(n18892) );
  INV_X1 U654 ( .A(n1142), .ZN(n18903) );
  NOR3_X1 U655 ( .A1(n3926), .A2(ADD_RD1[0]), .A3(n3928), .ZN(n3909) );
  NOR3_X1 U656 ( .A1(n3926), .A2(ADD_RD1[3]), .A3(n3929), .ZN(n3908) );
  NOR3_X1 U657 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(ADD_RD1[0]), .ZN(n3911)
         );
  NOR3_X1 U658 ( .A1(n3929), .A2(ADD_RD1[4]), .A3(n3928), .ZN(n3913) );
  NOR3_X1 U659 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(n3929), .ZN(n3915) );
  NOR3_X1 U660 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[3]), .A3(n3926), .ZN(n3912) );
  NOR3_X1 U661 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(n3928), .ZN(n3905) );
  INV_X1 U662 ( .A(n17839), .ZN(n18440) );
  INV_X1 U663 ( .A(n18352), .ZN(n18538) );
  OAI222_X1 U664 ( .A1(n18160), .A2(n18385), .B1(n17423), .B2(n18382), .C1(
        n17807), .C2(n18379), .ZN(n4102) );
  OAI222_X1 U665 ( .A1(n18161), .A2(n18385), .B1(n17424), .B2(n18382), .C1(
        n17808), .C2(n18379), .ZN(n4084) );
  OAI222_X1 U666 ( .A1(n18162), .A2(n18385), .B1(n17425), .B2(n18382), .C1(
        n17809), .C2(n18379), .ZN(n4066) );
  OAI222_X1 U667 ( .A1(n18163), .A2(n18385), .B1(n17426), .B2(n18382), .C1(
        n17810), .C2(n18379), .ZN(n4048) );
  OAI222_X1 U668 ( .A1(n18164), .A2(n18385), .B1(n17427), .B2(n18382), .C1(
        n17811), .C2(n18379), .ZN(n4030) );
  OAI222_X1 U669 ( .A1(n18165), .A2(n18385), .B1(n17428), .B2(n18382), .C1(
        n17812), .C2(n18379), .ZN(n4012) );
  OAI222_X1 U670 ( .A1(n18166), .A2(n18385), .B1(n17429), .B2(n18382), .C1(
        n17813), .C2(n18379), .ZN(n3994) );
  OAI222_X1 U671 ( .A1(n18167), .A2(n18385), .B1(n17430), .B2(n18382), .C1(
        n17814), .C2(n18379), .ZN(n3959) );
  OAI222_X1 U672 ( .A1(n18215), .A2(n18483), .B1(n17775), .B2(n18480), .C1(
        n17455), .C2(n18477), .ZN(n2364) );
  OAI222_X1 U673 ( .A1(n18216), .A2(n18483), .B1(n17776), .B2(n18480), .C1(
        n17456), .C2(n18477), .ZN(n2345) );
  OAI222_X1 U674 ( .A1(n18217), .A2(n18483), .B1(n17777), .B2(n18480), .C1(
        n17457), .C2(n18477), .ZN(n2326) );
  OAI222_X1 U675 ( .A1(n18218), .A2(n18483), .B1(n17778), .B2(n18480), .C1(
        n17458), .C2(n18477), .ZN(n2307) );
  OAI222_X1 U676 ( .A1(n18219), .A2(n18483), .B1(n17779), .B2(n18480), .C1(
        n17459), .C2(n18477), .ZN(n2288) );
  OAI222_X1 U677 ( .A1(n18220), .A2(n18483), .B1(n17780), .B2(n18480), .C1(
        n17460), .C2(n18477), .ZN(n2269) );
  OAI222_X1 U678 ( .A1(n18221), .A2(n18483), .B1(n17781), .B2(n18480), .C1(
        n17461), .C2(n18477), .ZN(n2250) );
  OAI222_X1 U679 ( .A1(n18222), .A2(n18483), .B1(n17782), .B2(n18480), .C1(
        n17462), .C2(n18477), .ZN(n2214) );
  OAI222_X1 U680 ( .A1(n18170), .A2(n18383), .B1(n17431), .B2(n18380), .C1(
        n17817), .C2(n18377), .ZN(n4546) );
  OAI222_X1 U681 ( .A1(n18168), .A2(n18383), .B1(n17433), .B2(n18380), .C1(
        n17818), .C2(n18377), .ZN(n4516) );
  OAI222_X1 U682 ( .A1(n18171), .A2(n18383), .B1(n17432), .B2(n18380), .C1(
        n17819), .C2(n18377), .ZN(n4498) );
  OAI222_X1 U683 ( .A1(n18172), .A2(n18383), .B1(n17434), .B2(n18380), .C1(
        n17815), .C2(n18377), .ZN(n4480) );
  OAI222_X1 U684 ( .A1(n18169), .A2(n18383), .B1(n17435), .B2(n18380), .C1(
        n17816), .C2(n18377), .ZN(n4462) );
  OAI222_X1 U685 ( .A1(n18173), .A2(n18383), .B1(n17436), .B2(n18380), .C1(
        n17820), .C2(n18377), .ZN(n4444) );
  OAI222_X1 U686 ( .A1(n18174), .A2(n18383), .B1(n17437), .B2(n18380), .C1(
        n17821), .C2(n18377), .ZN(n4426) );
  OAI222_X1 U687 ( .A1(n18175), .A2(n18383), .B1(n17438), .B2(n18380), .C1(
        n17822), .C2(n18377), .ZN(n4408) );
  OAI222_X1 U688 ( .A1(n18176), .A2(n18383), .B1(n17439), .B2(n18380), .C1(
        n17823), .C2(n18377), .ZN(n4390) );
  OAI222_X1 U689 ( .A1(n18177), .A2(n18383), .B1(n17440), .B2(n18380), .C1(
        n17824), .C2(n18377), .ZN(n4372) );
  OAI222_X1 U690 ( .A1(n18178), .A2(n18383), .B1(n17441), .B2(n18380), .C1(
        n17825), .C2(n18377), .ZN(n4354) );
  OAI222_X1 U691 ( .A1(n18179), .A2(n18383), .B1(n17442), .B2(n18380), .C1(
        n17826), .C2(n18377), .ZN(n4336) );
  OAI222_X1 U692 ( .A1(n18180), .A2(n18384), .B1(n17443), .B2(n18381), .C1(
        n17827), .C2(n18378), .ZN(n4318) );
  OAI222_X1 U693 ( .A1(n18181), .A2(n18384), .B1(n17444), .B2(n18381), .C1(
        n17828), .C2(n18378), .ZN(n4300) );
  OAI222_X1 U694 ( .A1(n18182), .A2(n18384), .B1(n17445), .B2(n18381), .C1(
        n17829), .C2(n18378), .ZN(n4282) );
  OAI222_X1 U695 ( .A1(n18183), .A2(n18384), .B1(n17446), .B2(n18381), .C1(
        n17830), .C2(n18378), .ZN(n4264) );
  OAI222_X1 U696 ( .A1(n18184), .A2(n18384), .B1(n17447), .B2(n18381), .C1(
        n17831), .C2(n18378), .ZN(n4246) );
  OAI222_X1 U697 ( .A1(n18185), .A2(n18384), .B1(n17448), .B2(n18381), .C1(
        n17832), .C2(n18378), .ZN(n4228) );
  OAI222_X1 U698 ( .A1(n18186), .A2(n18384), .B1(n17449), .B2(n18381), .C1(
        n17833), .C2(n18378), .ZN(n4210) );
  OAI222_X1 U699 ( .A1(n18187), .A2(n18384), .B1(n17450), .B2(n18381), .C1(
        n17834), .C2(n18378), .ZN(n4192) );
  OAI222_X1 U700 ( .A1(n18188), .A2(n18384), .B1(n17451), .B2(n18381), .C1(
        n17835), .C2(n18378), .ZN(n4174) );
  OAI222_X1 U701 ( .A1(n18189), .A2(n18384), .B1(n17452), .B2(n18381), .C1(
        n17836), .C2(n18378), .ZN(n4156) );
  OAI222_X1 U702 ( .A1(n18190), .A2(n18384), .B1(n17453), .B2(n18381), .C1(
        n17837), .C2(n18378), .ZN(n4138) );
  OAI222_X1 U703 ( .A1(n18191), .A2(n18384), .B1(n17454), .B2(n18381), .C1(
        n17838), .C2(n18378), .ZN(n4120) );
  OAI222_X1 U704 ( .A1(n18192), .A2(n18481), .B1(n17783), .B2(n18478), .C1(
        n17463), .C2(n18475), .ZN(n3920) );
  OAI222_X1 U705 ( .A1(n18193), .A2(n18481), .B1(n17785), .B2(n18478), .C1(
        n17467), .C2(n18475), .ZN(n3889) );
  OAI222_X1 U706 ( .A1(n18194), .A2(n18481), .B1(n17786), .B2(n18478), .C1(
        n17464), .C2(n18475), .ZN(n3870) );
  OAI222_X1 U707 ( .A1(n18286), .A2(n18481), .B1(n17784), .B2(n18478), .C1(
        n17465), .C2(n18475), .ZN(n3851) );
  OAI222_X1 U708 ( .A1(n18195), .A2(n18481), .B1(n17787), .B2(n18478), .C1(
        n17466), .C2(n18475), .ZN(n2744) );
  OAI222_X1 U709 ( .A1(n18196), .A2(n18481), .B1(n17788), .B2(n18478), .C1(
        n17468), .C2(n18475), .ZN(n2725) );
  OAI222_X1 U710 ( .A1(n18197), .A2(n18481), .B1(n17789), .B2(n18478), .C1(
        n17469), .C2(n18475), .ZN(n2706) );
  OAI222_X1 U711 ( .A1(n18198), .A2(n18481), .B1(n17790), .B2(n18478), .C1(
        n17470), .C2(n18475), .ZN(n2687) );
  OAI222_X1 U712 ( .A1(n18199), .A2(n18481), .B1(n17791), .B2(n18478), .C1(
        n17471), .C2(n18475), .ZN(n2668) );
  OAI222_X1 U713 ( .A1(n18200), .A2(n18481), .B1(n17792), .B2(n18478), .C1(
        n17472), .C2(n18475), .ZN(n2649) );
  OAI222_X1 U714 ( .A1(n18201), .A2(n18481), .B1(n17793), .B2(n18478), .C1(
        n17473), .C2(n18475), .ZN(n2630) );
  OAI222_X1 U715 ( .A1(n18202), .A2(n18481), .B1(n17794), .B2(n18478), .C1(
        n17474), .C2(n18475), .ZN(n2611) );
  OAI222_X1 U716 ( .A1(n18203), .A2(n18482), .B1(n17795), .B2(n18479), .C1(
        n17475), .C2(n18476), .ZN(n2592) );
  OAI222_X1 U717 ( .A1(n18204), .A2(n18482), .B1(n17796), .B2(n18479), .C1(
        n17476), .C2(n18476), .ZN(n2573) );
  OAI222_X1 U718 ( .A1(n18205), .A2(n18482), .B1(n17797), .B2(n18479), .C1(
        n17477), .C2(n18476), .ZN(n2554) );
  OAI222_X1 U719 ( .A1(n18206), .A2(n18482), .B1(n17798), .B2(n18479), .C1(
        n17478), .C2(n18476), .ZN(n2535) );
  OAI222_X1 U720 ( .A1(n18207), .A2(n18482), .B1(n17799), .B2(n18479), .C1(
        n17479), .C2(n18476), .ZN(n2516) );
  OAI222_X1 U721 ( .A1(n18208), .A2(n18482), .B1(n17800), .B2(n18479), .C1(
        n17480), .C2(n18476), .ZN(n2497) );
  OAI222_X1 U722 ( .A1(n18209), .A2(n18482), .B1(n17801), .B2(n18479), .C1(
        n17481), .C2(n18476), .ZN(n2478) );
  OAI222_X1 U723 ( .A1(n18210), .A2(n18482), .B1(n17802), .B2(n18479), .C1(
        n17482), .C2(n18476), .ZN(n2459) );
  OAI222_X1 U724 ( .A1(n18211), .A2(n18482), .B1(n17803), .B2(n18479), .C1(
        n17483), .C2(n18476), .ZN(n2440) );
  OAI222_X1 U725 ( .A1(n18212), .A2(n18482), .B1(n17804), .B2(n18479), .C1(
        n17484), .C2(n18476), .ZN(n2421) );
  OAI222_X1 U726 ( .A1(n18213), .A2(n18482), .B1(n17805), .B2(n18479), .C1(
        n17485), .C2(n18476), .ZN(n2402) );
  OAI222_X1 U727 ( .A1(n18214), .A2(n18482), .B1(n17806), .B2(n18479), .C1(
        n17486), .C2(n18476), .ZN(n2383) );
  NOR4_X1 U728 ( .A1(n4526), .A2(n4527), .A3(n4528), .A4(n4529), .ZN(n4525) );
  OAI221_X1 U729 ( .B1(n17463), .B2(n18437), .C1(n17535), .C2(n18434), .A(
        n4536), .ZN(n4528) );
  OAI221_X1 U730 ( .B1(n17402), .B2(n18425), .C1(n17638), .C2(n18422), .A(
        n4541), .ZN(n4527) );
  OAI221_X1 U731 ( .B1(n18138), .B2(n18448), .C1(n17583), .C2(n18445), .A(
        n4530), .ZN(n4529) );
  NOR4_X1 U732 ( .A1(n4508), .A2(n4509), .A3(n4510), .A4(n4511), .ZN(n4507) );
  OAI221_X1 U733 ( .B1(n17467), .B2(n18437), .C1(n17536), .C2(n18434), .A(
        n4513), .ZN(n4510) );
  OAI221_X1 U734 ( .B1(n17399), .B2(n18425), .C1(n17639), .C2(n18422), .A(
        n4514), .ZN(n4509) );
  OAI221_X1 U735 ( .B1(n18139), .B2(n18448), .C1(n17677), .C2(n18445), .A(
        n4512), .ZN(n4511) );
  NOR4_X1 U736 ( .A1(n4490), .A2(n4491), .A3(n4492), .A4(n4493), .ZN(n4489) );
  OAI221_X1 U737 ( .B1(n17464), .B2(n18437), .C1(n17540), .C2(n18434), .A(
        n4495), .ZN(n4492) );
  OAI221_X1 U738 ( .B1(n17400), .B2(n18425), .C1(n17678), .C2(n18422), .A(
        n4496), .ZN(n4491) );
  OAI221_X1 U739 ( .B1(n18136), .B2(n18448), .C1(n17584), .C2(n18445), .A(
        n4494), .ZN(n4493) );
  NOR4_X1 U740 ( .A1(n4472), .A2(n4473), .A3(n4474), .A4(n4475), .ZN(n4471) );
  OAI221_X1 U741 ( .B1(n17465), .B2(n18437), .C1(n17541), .C2(n18434), .A(
        n4477), .ZN(n4474) );
  OAI221_X1 U742 ( .B1(n17403), .B2(n18425), .C1(n17640), .C2(n18422), .A(
        n4478), .ZN(n4473) );
  OAI221_X1 U743 ( .B1(n18137), .B2(n18448), .C1(n17585), .C2(n18445), .A(
        n4476), .ZN(n4475) );
  NOR4_X1 U744 ( .A1(n4454), .A2(n4455), .A3(n4456), .A4(n4457), .ZN(n4453) );
  OAI221_X1 U745 ( .B1(n17466), .B2(n18437), .C1(n17542), .C2(n18434), .A(
        n4459), .ZN(n4456) );
  OAI221_X1 U746 ( .B1(n17401), .B2(n18425), .C1(n17641), .C2(n18422), .A(
        n4460), .ZN(n4455) );
  OAI221_X1 U747 ( .B1(n18140), .B2(n18448), .C1(n17586), .C2(n18445), .A(
        n4458), .ZN(n4457) );
  NOR4_X1 U748 ( .A1(n4436), .A2(n4437), .A3(n4438), .A4(n4439), .ZN(n4435) );
  OAI221_X1 U749 ( .B1(n17468), .B2(n18437), .C1(n17543), .C2(n18434), .A(
        n4441), .ZN(n4438) );
  OAI221_X1 U750 ( .B1(n17404), .B2(n18425), .C1(n17642), .C2(n18422), .A(
        n4442), .ZN(n4437) );
  OAI221_X1 U751 ( .B1(n18141), .B2(n18448), .C1(n17587), .C2(n18445), .A(
        n4440), .ZN(n4439) );
  NOR4_X1 U752 ( .A1(n4418), .A2(n4419), .A3(n4420), .A4(n4421), .ZN(n4417) );
  OAI221_X1 U753 ( .B1(n17469), .B2(n18437), .C1(n17544), .C2(n18434), .A(
        n4423), .ZN(n4420) );
  OAI221_X1 U754 ( .B1(n17405), .B2(n18425), .C1(n17643), .C2(n18422), .A(
        n4424), .ZN(n4419) );
  OAI221_X1 U755 ( .B1(n18142), .B2(n18448), .C1(n17588), .C2(n18445), .A(
        n4422), .ZN(n4421) );
  NOR4_X1 U756 ( .A1(n4400), .A2(n4401), .A3(n4402), .A4(n4403), .ZN(n4399) );
  OAI221_X1 U757 ( .B1(n17470), .B2(n18437), .C1(n17545), .C2(n18434), .A(
        n4405), .ZN(n4402) );
  OAI221_X1 U758 ( .B1(n17406), .B2(n18425), .C1(n17644), .C2(n18422), .A(
        n4406), .ZN(n4401) );
  OAI221_X1 U759 ( .B1(n18143), .B2(n18448), .C1(n17589), .C2(n18445), .A(
        n4404), .ZN(n4403) );
  NOR4_X1 U760 ( .A1(n4382), .A2(n4383), .A3(n4384), .A4(n4385), .ZN(n4381) );
  OAI221_X1 U761 ( .B1(n17471), .B2(n18437), .C1(n17546), .C2(n18434), .A(
        n4387), .ZN(n4384) );
  OAI221_X1 U762 ( .B1(n17407), .B2(n18425), .C1(n17645), .C2(n18422), .A(
        n4388), .ZN(n4383) );
  OAI221_X1 U763 ( .B1(n18144), .B2(n18448), .C1(n17590), .C2(n18445), .A(
        n4386), .ZN(n4385) );
  NOR4_X1 U764 ( .A1(n4364), .A2(n4365), .A3(n4366), .A4(n4367), .ZN(n4363) );
  OAI221_X1 U765 ( .B1(n17472), .B2(n18437), .C1(n17547), .C2(n18434), .A(
        n4369), .ZN(n4366) );
  OAI221_X1 U766 ( .B1(n17408), .B2(n18425), .C1(n17646), .C2(n18422), .A(
        n4370), .ZN(n4365) );
  OAI221_X1 U767 ( .B1(n18145), .B2(n18448), .C1(n17591), .C2(n18445), .A(
        n4368), .ZN(n4367) );
  NOR4_X1 U768 ( .A1(n4346), .A2(n4347), .A3(n4348), .A4(n4349), .ZN(n4345) );
  OAI221_X1 U769 ( .B1(n17473), .B2(n18437), .C1(n17548), .C2(n18434), .A(
        n4351), .ZN(n4348) );
  OAI221_X1 U770 ( .B1(n17409), .B2(n18425), .C1(n17647), .C2(n18422), .A(
        n4352), .ZN(n4347) );
  OAI221_X1 U771 ( .B1(n18146), .B2(n18448), .C1(n17592), .C2(n18445), .A(
        n4350), .ZN(n4349) );
  NOR4_X1 U772 ( .A1(n4328), .A2(n4329), .A3(n4330), .A4(n4331), .ZN(n4327) );
  OAI221_X1 U773 ( .B1(n17474), .B2(n18437), .C1(n17549), .C2(n18434), .A(
        n4333), .ZN(n4330) );
  OAI221_X1 U774 ( .B1(n17410), .B2(n18425), .C1(n17648), .C2(n18422), .A(
        n4334), .ZN(n4329) );
  OAI221_X1 U775 ( .B1(n18147), .B2(n18448), .C1(n17593), .C2(n18445), .A(
        n4332), .ZN(n4331) );
  NOR4_X1 U776 ( .A1(n4310), .A2(n4311), .A3(n4312), .A4(n4313), .ZN(n4309) );
  OAI221_X1 U777 ( .B1(n17475), .B2(n18438), .C1(n17550), .C2(n18435), .A(
        n4315), .ZN(n4312) );
  OAI221_X1 U778 ( .B1(n17411), .B2(n18426), .C1(n17649), .C2(n18423), .A(
        n4316), .ZN(n4311) );
  OAI221_X1 U779 ( .B1(n18148), .B2(n18449), .C1(n17594), .C2(n18446), .A(
        n4314), .ZN(n4313) );
  NOR4_X1 U780 ( .A1(n4292), .A2(n4293), .A3(n4294), .A4(n4295), .ZN(n4291) );
  OAI221_X1 U781 ( .B1(n17476), .B2(n18438), .C1(n17551), .C2(n18435), .A(
        n4297), .ZN(n4294) );
  OAI221_X1 U782 ( .B1(n17412), .B2(n18426), .C1(n17650), .C2(n18423), .A(
        n4298), .ZN(n4293) );
  OAI221_X1 U783 ( .B1(n18149), .B2(n18449), .C1(n17595), .C2(n18446), .A(
        n4296), .ZN(n4295) );
  NOR4_X1 U784 ( .A1(n4274), .A2(n4275), .A3(n4276), .A4(n4277), .ZN(n4273) );
  OAI221_X1 U785 ( .B1(n17477), .B2(n18438), .C1(n17552), .C2(n18435), .A(
        n4279), .ZN(n4276) );
  OAI221_X1 U786 ( .B1(n17413), .B2(n18426), .C1(n17651), .C2(n18423), .A(
        n4280), .ZN(n4275) );
  OAI221_X1 U787 ( .B1(n18150), .B2(n18449), .C1(n17596), .C2(n18446), .A(
        n4278), .ZN(n4277) );
  NOR4_X1 U788 ( .A1(n4256), .A2(n4257), .A3(n4258), .A4(n4259), .ZN(n4255) );
  OAI221_X1 U789 ( .B1(n17478), .B2(n18438), .C1(n17553), .C2(n18435), .A(
        n4261), .ZN(n4258) );
  OAI221_X1 U790 ( .B1(n17414), .B2(n18426), .C1(n17652), .C2(n18423), .A(
        n4262), .ZN(n4257) );
  OAI221_X1 U791 ( .B1(n18151), .B2(n18449), .C1(n17597), .C2(n18446), .A(
        n4260), .ZN(n4259) );
  NOR4_X1 U792 ( .A1(n4238), .A2(n4239), .A3(n4240), .A4(n4241), .ZN(n4237) );
  OAI221_X1 U793 ( .B1(n17479), .B2(n18438), .C1(n17554), .C2(n18435), .A(
        n4243), .ZN(n4240) );
  OAI221_X1 U794 ( .B1(n17415), .B2(n18426), .C1(n17653), .C2(n18423), .A(
        n4244), .ZN(n4239) );
  OAI221_X1 U795 ( .B1(n18152), .B2(n18449), .C1(n17598), .C2(n18446), .A(
        n4242), .ZN(n4241) );
  NOR4_X1 U796 ( .A1(n4220), .A2(n4221), .A3(n4222), .A4(n4223), .ZN(n4219) );
  OAI221_X1 U797 ( .B1(n17480), .B2(n18438), .C1(n17555), .C2(n18435), .A(
        n4225), .ZN(n4222) );
  OAI221_X1 U798 ( .B1(n17416), .B2(n18426), .C1(n17654), .C2(n18423), .A(
        n4226), .ZN(n4221) );
  OAI221_X1 U799 ( .B1(n18153), .B2(n18449), .C1(n17599), .C2(n18446), .A(
        n4224), .ZN(n4223) );
  NOR4_X1 U800 ( .A1(n4202), .A2(n4203), .A3(n4204), .A4(n4205), .ZN(n4201) );
  OAI221_X1 U801 ( .B1(n17481), .B2(n18438), .C1(n17556), .C2(n18435), .A(
        n4207), .ZN(n4204) );
  OAI221_X1 U802 ( .B1(n17417), .B2(n18426), .C1(n17655), .C2(n18423), .A(
        n4208), .ZN(n4203) );
  OAI221_X1 U803 ( .B1(n18154), .B2(n18449), .C1(n17600), .C2(n18446), .A(
        n4206), .ZN(n4205) );
  NOR4_X1 U804 ( .A1(n4184), .A2(n4185), .A3(n4186), .A4(n4187), .ZN(n4183) );
  OAI221_X1 U805 ( .B1(n17482), .B2(n18438), .C1(n17557), .C2(n18435), .A(
        n4189), .ZN(n4186) );
  OAI221_X1 U806 ( .B1(n17418), .B2(n18426), .C1(n17656), .C2(n18423), .A(
        n4190), .ZN(n4185) );
  OAI221_X1 U807 ( .B1(n18155), .B2(n18449), .C1(n17601), .C2(n18446), .A(
        n4188), .ZN(n4187) );
  NOR4_X1 U808 ( .A1(n4166), .A2(n4167), .A3(n4168), .A4(n4169), .ZN(n4165) );
  OAI221_X1 U809 ( .B1(n17483), .B2(n18438), .C1(n17558), .C2(n18435), .A(
        n4171), .ZN(n4168) );
  OAI221_X1 U810 ( .B1(n17419), .B2(n18426), .C1(n17657), .C2(n18423), .A(
        n4172), .ZN(n4167) );
  OAI221_X1 U811 ( .B1(n18156), .B2(n18449), .C1(n17602), .C2(n18446), .A(
        n4170), .ZN(n4169) );
  NOR4_X1 U812 ( .A1(n4148), .A2(n4149), .A3(n4150), .A4(n4151), .ZN(n4147) );
  OAI221_X1 U813 ( .B1(n17484), .B2(n18438), .C1(n17559), .C2(n18435), .A(
        n4153), .ZN(n4150) );
  OAI221_X1 U814 ( .B1(n17420), .B2(n18426), .C1(n17658), .C2(n18423), .A(
        n4154), .ZN(n4149) );
  OAI221_X1 U815 ( .B1(n18157), .B2(n18449), .C1(n17603), .C2(n18446), .A(
        n4152), .ZN(n4151) );
  NOR4_X1 U816 ( .A1(n4130), .A2(n4131), .A3(n4132), .A4(n4133), .ZN(n4129) );
  OAI221_X1 U817 ( .B1(n17485), .B2(n18438), .C1(n17560), .C2(n18435), .A(
        n4135), .ZN(n4132) );
  OAI221_X1 U818 ( .B1(n17421), .B2(n18426), .C1(n17659), .C2(n18423), .A(
        n4136), .ZN(n4131) );
  OAI221_X1 U819 ( .B1(n18158), .B2(n18449), .C1(n17604), .C2(n18446), .A(
        n4134), .ZN(n4133) );
  NOR4_X1 U820 ( .A1(n4112), .A2(n4113), .A3(n4114), .A4(n4115), .ZN(n4111) );
  OAI221_X1 U821 ( .B1(n17486), .B2(n18438), .C1(n17561), .C2(n18435), .A(
        n4117), .ZN(n4114) );
  OAI221_X1 U822 ( .B1(n17422), .B2(n18426), .C1(n17660), .C2(n18423), .A(
        n4118), .ZN(n4113) );
  OAI221_X1 U823 ( .B1(n18159), .B2(n18449), .C1(n17605), .C2(n18446), .A(
        n4116), .ZN(n4115) );
  NOR4_X1 U824 ( .A1(n3900), .A2(n3901), .A3(n3902), .A4(n3903), .ZN(n3899) );
  OAI221_X1 U825 ( .B1(n17754), .B2(n18511), .C1(n18262), .C2(n18508), .A(
        n3918), .ZN(n3900) );
  OAI221_X1 U826 ( .B1(n17431), .B2(n18523), .C1(n17537), .C2(n18520), .A(
        n3916), .ZN(n3901) );
  OAI221_X1 U827 ( .B1(n17715), .B2(n18535), .C1(n18223), .C2(n18532), .A(
        n3910), .ZN(n3902) );
  NOR4_X1 U828 ( .A1(n3881), .A2(n3882), .A3(n3883), .A4(n3884), .ZN(n3880) );
  OAI221_X1 U829 ( .B1(n17751), .B2(n18511), .C1(n18263), .C2(n18508), .A(
        n3888), .ZN(n3881) );
  OAI221_X1 U830 ( .B1(n17433), .B2(n18523), .C1(n17562), .C2(n18520), .A(
        n3887), .ZN(n3882) );
  OAI221_X1 U831 ( .B1(n17711), .B2(n18535), .C1(n18224), .C2(n18532), .A(
        n3886), .ZN(n3883) );
  NOR4_X1 U832 ( .A1(n3862), .A2(n3863), .A3(n3864), .A4(n3865), .ZN(n3861) );
  OAI221_X1 U833 ( .B1(n17752), .B2(n18511), .C1(n18266), .C2(n18508), .A(
        n3869), .ZN(n3862) );
  OAI221_X1 U834 ( .B1(n17432), .B2(n18523), .C1(n17538), .C2(n18520), .A(
        n3868), .ZN(n3863) );
  OAI221_X1 U835 ( .B1(n17712), .B2(n18535), .C1(n18225), .C2(n18532), .A(
        n3867), .ZN(n3864) );
  NOR4_X1 U836 ( .A1(n2755), .A2(n2756), .A3(n2757), .A4(n2758), .ZN(n2754) );
  OAI221_X1 U837 ( .B1(n17753), .B2(n18511), .C1(n18264), .C2(n18508), .A(
        n3850), .ZN(n2755) );
  OAI221_X1 U838 ( .B1(n17434), .B2(n18523), .C1(n17563), .C2(n18520), .A(
        n3849), .ZN(n2756) );
  OAI221_X1 U839 ( .B1(n17713), .B2(n18535), .C1(n18226), .C2(n18532), .A(
        n3848), .ZN(n2757) );
  NOR4_X1 U840 ( .A1(n2736), .A2(n2737), .A3(n2738), .A4(n2739), .ZN(n2735) );
  OAI221_X1 U841 ( .B1(n17755), .B2(n18511), .C1(n18265), .C2(n18508), .A(
        n2743), .ZN(n2736) );
  OAI221_X1 U842 ( .B1(n17435), .B2(n18523), .C1(n17539), .C2(n18520), .A(
        n2742), .ZN(n2737) );
  OAI221_X1 U843 ( .B1(n17714), .B2(n18535), .C1(n18287), .C2(n18532), .A(
        n2741), .ZN(n2738) );
  NOR4_X1 U844 ( .A1(n2717), .A2(n2718), .A3(n2719), .A4(n2720), .ZN(n2716) );
  OAI221_X1 U845 ( .B1(n17756), .B2(n18511), .C1(n18267), .C2(n18508), .A(
        n2724), .ZN(n2717) );
  OAI221_X1 U846 ( .B1(n17436), .B2(n18523), .C1(n17564), .C2(n18520), .A(
        n2723), .ZN(n2718) );
  OAI221_X1 U847 ( .B1(n17716), .B2(n18535), .C1(n18227), .C2(n18532), .A(
        n2722), .ZN(n2719) );
  NOR4_X1 U848 ( .A1(n2698), .A2(n2699), .A3(n2700), .A4(n2701), .ZN(n2697) );
  OAI221_X1 U849 ( .B1(n17757), .B2(n18511), .C1(n18268), .C2(n18508), .A(
        n2705), .ZN(n2698) );
  OAI221_X1 U850 ( .B1(n17437), .B2(n18523), .C1(n17565), .C2(n18520), .A(
        n2704), .ZN(n2699) );
  OAI221_X1 U851 ( .B1(n17717), .B2(n18535), .C1(n18228), .C2(n18532), .A(
        n2703), .ZN(n2700) );
  NOR4_X1 U852 ( .A1(n2679), .A2(n2680), .A3(n2681), .A4(n2682), .ZN(n2678) );
  OAI221_X1 U853 ( .B1(n17758), .B2(n18511), .C1(n18269), .C2(n18508), .A(
        n2686), .ZN(n2679) );
  OAI221_X1 U854 ( .B1(n17438), .B2(n18523), .C1(n17566), .C2(n18520), .A(
        n2685), .ZN(n2680) );
  OAI221_X1 U855 ( .B1(n17718), .B2(n18535), .C1(n18229), .C2(n18532), .A(
        n2684), .ZN(n2681) );
  NOR4_X1 U856 ( .A1(n2660), .A2(n2661), .A3(n2662), .A4(n2663), .ZN(n2659) );
  OAI221_X1 U857 ( .B1(n17759), .B2(n18511), .C1(n18270), .C2(n18508), .A(
        n2667), .ZN(n2660) );
  OAI221_X1 U858 ( .B1(n17439), .B2(n18523), .C1(n17567), .C2(n18520), .A(
        n2666), .ZN(n2661) );
  OAI221_X1 U859 ( .B1(n17367), .B2(n18546), .C1(n17622), .C2(n18543), .A(
        n2664), .ZN(n2663) );
  NOR4_X1 U860 ( .A1(n2641), .A2(n2642), .A3(n2643), .A4(n2644), .ZN(n2640) );
  OAI221_X1 U861 ( .B1(n17760), .B2(n18511), .C1(n18271), .C2(n18508), .A(
        n2648), .ZN(n2641) );
  OAI221_X1 U862 ( .B1(n17440), .B2(n18523), .C1(n17568), .C2(n18520), .A(
        n2647), .ZN(n2642) );
  OAI221_X1 U863 ( .B1(n17368), .B2(n18546), .C1(n17623), .C2(n18543), .A(
        n2645), .ZN(n2644) );
  NOR4_X1 U864 ( .A1(n2622), .A2(n2623), .A3(n2624), .A4(n2625), .ZN(n2621) );
  OAI221_X1 U865 ( .B1(n17761), .B2(n18511), .C1(n18272), .C2(n18508), .A(
        n2629), .ZN(n2622) );
  OAI221_X1 U866 ( .B1(n17441), .B2(n18523), .C1(n17569), .C2(n18520), .A(
        n2628), .ZN(n2623) );
  OAI221_X1 U867 ( .B1(n17369), .B2(n18546), .C1(n17624), .C2(n18543), .A(
        n2626), .ZN(n2625) );
  NOR4_X1 U868 ( .A1(n2603), .A2(n2604), .A3(n2605), .A4(n2606), .ZN(n2602) );
  OAI221_X1 U869 ( .B1(n17762), .B2(n18511), .C1(n18273), .C2(n18508), .A(
        n2610), .ZN(n2603) );
  OAI221_X1 U870 ( .B1(n17442), .B2(n18523), .C1(n17570), .C2(n18520), .A(
        n2609), .ZN(n2604) );
  OAI221_X1 U871 ( .B1(n17370), .B2(n18546), .C1(n17625), .C2(n18543), .A(
        n2607), .ZN(n2606) );
  NOR4_X1 U872 ( .A1(n2584), .A2(n2585), .A3(n2586), .A4(n2587), .ZN(n2583) );
  OAI221_X1 U873 ( .B1(n17763), .B2(n18512), .C1(n18274), .C2(n18509), .A(
        n2591), .ZN(n2584) );
  OAI221_X1 U874 ( .B1(n17443), .B2(n18524), .C1(n17571), .C2(n18521), .A(
        n2590), .ZN(n2585) );
  OAI221_X1 U875 ( .B1(n17371), .B2(n18547), .C1(n17626), .C2(n18544), .A(
        n2588), .ZN(n2587) );
  NOR4_X1 U876 ( .A1(n2565), .A2(n2566), .A3(n2567), .A4(n2568), .ZN(n2564) );
  OAI221_X1 U877 ( .B1(n17764), .B2(n18512), .C1(n18275), .C2(n18509), .A(
        n2572), .ZN(n2565) );
  OAI221_X1 U878 ( .B1(n17444), .B2(n18524), .C1(n17572), .C2(n18521), .A(
        n2571), .ZN(n2566) );
  OAI221_X1 U879 ( .B1(n17372), .B2(n18547), .C1(n17627), .C2(n18544), .A(
        n2569), .ZN(n2568) );
  NOR4_X1 U880 ( .A1(n2546), .A2(n2547), .A3(n2548), .A4(n2549), .ZN(n2545) );
  OAI221_X1 U881 ( .B1(n17765), .B2(n18512), .C1(n18276), .C2(n18509), .A(
        n2553), .ZN(n2546) );
  OAI221_X1 U882 ( .B1(n17445), .B2(n18524), .C1(n17573), .C2(n18521), .A(
        n2552), .ZN(n2547) );
  OAI221_X1 U883 ( .B1(n17373), .B2(n18547), .C1(n17628), .C2(n18544), .A(
        n2550), .ZN(n2549) );
  NOR4_X1 U884 ( .A1(n2527), .A2(n2528), .A3(n2529), .A4(n2530), .ZN(n2526) );
  OAI221_X1 U885 ( .B1(n17766), .B2(n18512), .C1(n18277), .C2(n18509), .A(
        n2534), .ZN(n2527) );
  OAI221_X1 U886 ( .B1(n17446), .B2(n18524), .C1(n17574), .C2(n18521), .A(
        n2533), .ZN(n2528) );
  OAI221_X1 U887 ( .B1(n17374), .B2(n18547), .C1(n17629), .C2(n18544), .A(
        n2531), .ZN(n2530) );
  NOR4_X1 U888 ( .A1(n2508), .A2(n2509), .A3(n2510), .A4(n2511), .ZN(n2507) );
  OAI221_X1 U889 ( .B1(n17767), .B2(n18512), .C1(n18278), .C2(n18509), .A(
        n2515), .ZN(n2508) );
  OAI221_X1 U890 ( .B1(n17447), .B2(n18524), .C1(n17575), .C2(n18521), .A(
        n2514), .ZN(n2509) );
  OAI221_X1 U891 ( .B1(n17375), .B2(n18547), .C1(n17630), .C2(n18544), .A(
        n2512), .ZN(n2511) );
  NOR4_X1 U892 ( .A1(n2489), .A2(n2490), .A3(n2491), .A4(n2492), .ZN(n2488) );
  OAI221_X1 U893 ( .B1(n17768), .B2(n18512), .C1(n18279), .C2(n18509), .A(
        n2496), .ZN(n2489) );
  OAI221_X1 U894 ( .B1(n17448), .B2(n18524), .C1(n17576), .C2(n18521), .A(
        n2495), .ZN(n2490) );
  OAI221_X1 U895 ( .B1(n17376), .B2(n18547), .C1(n17631), .C2(n18544), .A(
        n2493), .ZN(n2492) );
  NOR4_X1 U896 ( .A1(n2470), .A2(n2471), .A3(n2472), .A4(n2473), .ZN(n2469) );
  OAI221_X1 U897 ( .B1(n17769), .B2(n18512), .C1(n18280), .C2(n18509), .A(
        n2477), .ZN(n2470) );
  OAI221_X1 U898 ( .B1(n17449), .B2(n18524), .C1(n17577), .C2(n18521), .A(
        n2476), .ZN(n2471) );
  OAI221_X1 U899 ( .B1(n17377), .B2(n18547), .C1(n17632), .C2(n18544), .A(
        n2474), .ZN(n2473) );
  NOR4_X1 U900 ( .A1(n2451), .A2(n2452), .A3(n2453), .A4(n2454), .ZN(n2450) );
  OAI221_X1 U901 ( .B1(n17770), .B2(n18512), .C1(n18281), .C2(n18509), .A(
        n2458), .ZN(n2451) );
  OAI221_X1 U902 ( .B1(n17450), .B2(n18524), .C1(n17578), .C2(n18521), .A(
        n2457), .ZN(n2452) );
  OAI221_X1 U903 ( .B1(n17378), .B2(n18547), .C1(n17633), .C2(n18544), .A(
        n2455), .ZN(n2454) );
  NOR4_X1 U904 ( .A1(n2432), .A2(n2433), .A3(n2434), .A4(n2435), .ZN(n2431) );
  OAI221_X1 U905 ( .B1(n17771), .B2(n18512), .C1(n18282), .C2(n18509), .A(
        n2439), .ZN(n2432) );
  OAI221_X1 U906 ( .B1(n17451), .B2(n18524), .C1(n17579), .C2(n18521), .A(
        n2438), .ZN(n2433) );
  OAI221_X1 U907 ( .B1(n17379), .B2(n18547), .C1(n17634), .C2(n18544), .A(
        n2436), .ZN(n2435) );
  NOR4_X1 U908 ( .A1(n2413), .A2(n2414), .A3(n2415), .A4(n2416), .ZN(n2412) );
  OAI221_X1 U909 ( .B1(n17772), .B2(n18512), .C1(n18283), .C2(n18509), .A(
        n2420), .ZN(n2413) );
  OAI221_X1 U910 ( .B1(n17452), .B2(n18524), .C1(n17580), .C2(n18521), .A(
        n2419), .ZN(n2414) );
  OAI221_X1 U911 ( .B1(n17380), .B2(n18547), .C1(n17635), .C2(n18544), .A(
        n2417), .ZN(n2416) );
  NOR4_X1 U912 ( .A1(n2394), .A2(n2395), .A3(n2396), .A4(n2397), .ZN(n2393) );
  OAI221_X1 U913 ( .B1(n17773), .B2(n18512), .C1(n18284), .C2(n18509), .A(
        n2401), .ZN(n2394) );
  OAI221_X1 U914 ( .B1(n17453), .B2(n18524), .C1(n17581), .C2(n18521), .A(
        n2400), .ZN(n2395) );
  OAI221_X1 U915 ( .B1(n17381), .B2(n18547), .C1(n17636), .C2(n18544), .A(
        n2398), .ZN(n2397) );
  NOR4_X1 U916 ( .A1(n2375), .A2(n2376), .A3(n2377), .A4(n2378), .ZN(n2374) );
  OAI221_X1 U917 ( .B1(n17774), .B2(n18512), .C1(n18285), .C2(n18509), .A(
        n2382), .ZN(n2375) );
  OAI221_X1 U918 ( .B1(n17454), .B2(n18524), .C1(n17582), .C2(n18521), .A(
        n2381), .ZN(n2376) );
  OAI221_X1 U919 ( .B1(n17382), .B2(n18547), .C1(n17637), .C2(n18544), .A(
        n2379), .ZN(n2378) );
  NOR4_X1 U920 ( .A1(n4094), .A2(n4095), .A3(n4096), .A4(n4097), .ZN(n4093) );
  OAI221_X1 U921 ( .B1(n17455), .B2(n18439), .C1(n17519), .C2(n18436), .A(
        n4099), .ZN(n4096) );
  OAI221_X1 U922 ( .B1(n18128), .B2(n18450), .C1(n17606), .C2(n18447), .A(
        n4098), .ZN(n4097) );
  OAI221_X1 U923 ( .B1(n17391), .B2(n18427), .C1(n17661), .C2(n18424), .A(
        n4100), .ZN(n4095) );
  NOR4_X1 U924 ( .A1(n4076), .A2(n4077), .A3(n4078), .A4(n4079), .ZN(n4075) );
  OAI221_X1 U925 ( .B1(n17456), .B2(n18439), .C1(n17520), .C2(n18436), .A(
        n4081), .ZN(n4078) );
  OAI221_X1 U926 ( .B1(n18129), .B2(n18450), .C1(n17607), .C2(n18447), .A(
        n4080), .ZN(n4079) );
  OAI221_X1 U927 ( .B1(n17392), .B2(n18427), .C1(n17662), .C2(n18424), .A(
        n4082), .ZN(n4077) );
  NOR4_X1 U928 ( .A1(n4058), .A2(n4059), .A3(n4060), .A4(n4061), .ZN(n4057) );
  OAI221_X1 U929 ( .B1(n17457), .B2(n18439), .C1(n17521), .C2(n18436), .A(
        n4063), .ZN(n4060) );
  OAI221_X1 U930 ( .B1(n18130), .B2(n18450), .C1(n17608), .C2(n18447), .A(
        n4062), .ZN(n4061) );
  OAI221_X1 U931 ( .B1(n17393), .B2(n18427), .C1(n17663), .C2(n18424), .A(
        n4064), .ZN(n4059) );
  NOR4_X1 U932 ( .A1(n4040), .A2(n4041), .A3(n4042), .A4(n4043), .ZN(n4039) );
  OAI221_X1 U933 ( .B1(n17458), .B2(n18439), .C1(n17522), .C2(n18436), .A(
        n4045), .ZN(n4042) );
  OAI221_X1 U934 ( .B1(n18131), .B2(n18450), .C1(n17609), .C2(n18447), .A(
        n4044), .ZN(n4043) );
  OAI221_X1 U935 ( .B1(n17394), .B2(n18427), .C1(n17664), .C2(n18424), .A(
        n4046), .ZN(n4041) );
  NOR4_X1 U936 ( .A1(n4022), .A2(n4023), .A3(n4024), .A4(n4025), .ZN(n4021) );
  OAI221_X1 U937 ( .B1(n17459), .B2(n18439), .C1(n17523), .C2(n18436), .A(
        n4027), .ZN(n4024) );
  OAI221_X1 U938 ( .B1(n18132), .B2(n18450), .C1(n17610), .C2(n18447), .A(
        n4026), .ZN(n4025) );
  OAI221_X1 U939 ( .B1(n17395), .B2(n18427), .C1(n17665), .C2(n18424), .A(
        n4028), .ZN(n4023) );
  NOR4_X1 U940 ( .A1(n4004), .A2(n4005), .A3(n4006), .A4(n4007), .ZN(n4003) );
  OAI221_X1 U941 ( .B1(n17460), .B2(n18439), .C1(n17524), .C2(n18436), .A(
        n4009), .ZN(n4006) );
  OAI221_X1 U942 ( .B1(n18133), .B2(n18450), .C1(n17611), .C2(n18447), .A(
        n4008), .ZN(n4007) );
  OAI221_X1 U943 ( .B1(n17396), .B2(n18427), .C1(n17666), .C2(n18424), .A(
        n4010), .ZN(n4005) );
  NOR4_X1 U944 ( .A1(n3986), .A2(n3987), .A3(n3988), .A4(n3989), .ZN(n3985) );
  OAI221_X1 U945 ( .B1(n17461), .B2(n18439), .C1(n17525), .C2(n18436), .A(
        n3991), .ZN(n3988) );
  OAI221_X1 U946 ( .B1(n18134), .B2(n18450), .C1(n17612), .C2(n18447), .A(
        n3990), .ZN(n3989) );
  OAI221_X1 U947 ( .B1(n17397), .B2(n18427), .C1(n17667), .C2(n18424), .A(
        n3992), .ZN(n3987) );
  NOR4_X1 U948 ( .A1(n3935), .A2(n3936), .A3(n3937), .A4(n3938), .ZN(n3934) );
  OAI221_X1 U949 ( .B1(n17462), .B2(n18439), .C1(n17526), .C2(n18436), .A(
        n3946), .ZN(n3937) );
  OAI221_X1 U950 ( .B1(n18135), .B2(n18450), .C1(n17613), .C2(n18447), .A(
        n3941), .ZN(n3938) );
  OAI221_X1 U951 ( .B1(n17398), .B2(n18427), .C1(n17668), .C2(n18424), .A(
        n3951), .ZN(n3936) );
  NOR4_X1 U952 ( .A1(n2356), .A2(n2357), .A3(n2358), .A4(n2359), .ZN(n2355) );
  OAI221_X1 U953 ( .B1(n17743), .B2(n18513), .C1(n18254), .C2(n18510), .A(
        n2363), .ZN(n2356) );
  OAI221_X1 U954 ( .B1(n17359), .B2(n18548), .C1(n17614), .C2(n18545), .A(
        n2360), .ZN(n2359) );
  OAI221_X1 U955 ( .B1(n17423), .B2(n18525), .C1(n17527), .C2(n18522), .A(
        n2362), .ZN(n2357) );
  NOR4_X1 U956 ( .A1(n2337), .A2(n2338), .A3(n2339), .A4(n2340), .ZN(n2336) );
  OAI221_X1 U957 ( .B1(n17744), .B2(n18513), .C1(n18255), .C2(n18510), .A(
        n2344), .ZN(n2337) );
  OAI221_X1 U958 ( .B1(n17360), .B2(n18548), .C1(n17615), .C2(n18545), .A(
        n2341), .ZN(n2340) );
  OAI221_X1 U959 ( .B1(n17424), .B2(n18525), .C1(n17528), .C2(n18522), .A(
        n2343), .ZN(n2338) );
  NOR4_X1 U960 ( .A1(n2318), .A2(n2319), .A3(n2320), .A4(n2321), .ZN(n2317) );
  OAI221_X1 U961 ( .B1(n17745), .B2(n18513), .C1(n18256), .C2(n18510), .A(
        n2325), .ZN(n2318) );
  OAI221_X1 U962 ( .B1(n17361), .B2(n18548), .C1(n17616), .C2(n18545), .A(
        n2322), .ZN(n2321) );
  OAI221_X1 U963 ( .B1(n17425), .B2(n18525), .C1(n17529), .C2(n18522), .A(
        n2324), .ZN(n2319) );
  NOR4_X1 U964 ( .A1(n2299), .A2(n2300), .A3(n2301), .A4(n2302), .ZN(n2298) );
  OAI221_X1 U965 ( .B1(n17746), .B2(n18513), .C1(n18257), .C2(n18510), .A(
        n2306), .ZN(n2299) );
  OAI221_X1 U966 ( .B1(n17362), .B2(n18548), .C1(n17617), .C2(n18545), .A(
        n2303), .ZN(n2302) );
  OAI221_X1 U967 ( .B1(n17426), .B2(n18525), .C1(n17530), .C2(n18522), .A(
        n2305), .ZN(n2300) );
  NOR4_X1 U968 ( .A1(n2280), .A2(n2281), .A3(n2282), .A4(n2283), .ZN(n2279) );
  OAI221_X1 U969 ( .B1(n17747), .B2(n18513), .C1(n18258), .C2(n18510), .A(
        n2287), .ZN(n2280) );
  OAI221_X1 U970 ( .B1(n17363), .B2(n18548), .C1(n17618), .C2(n18545), .A(
        n2284), .ZN(n2283) );
  OAI221_X1 U971 ( .B1(n17427), .B2(n18525), .C1(n17531), .C2(n18522), .A(
        n2286), .ZN(n2281) );
  NOR4_X1 U972 ( .A1(n2261), .A2(n2262), .A3(n2263), .A4(n2264), .ZN(n2260) );
  OAI221_X1 U973 ( .B1(n17748), .B2(n18513), .C1(n18259), .C2(n18510), .A(
        n2268), .ZN(n2261) );
  OAI221_X1 U974 ( .B1(n17364), .B2(n18548), .C1(n17619), .C2(n18545), .A(
        n2265), .ZN(n2264) );
  OAI221_X1 U975 ( .B1(n17428), .B2(n18525), .C1(n17532), .C2(n18522), .A(
        n2267), .ZN(n2262) );
  NOR4_X1 U976 ( .A1(n2242), .A2(n2243), .A3(n2244), .A4(n2245), .ZN(n2241) );
  OAI221_X1 U977 ( .B1(n17749), .B2(n18513), .C1(n18260), .C2(n18510), .A(
        n2249), .ZN(n2242) );
  OAI221_X1 U978 ( .B1(n17365), .B2(n18548), .C1(n17620), .C2(n18545), .A(
        n2246), .ZN(n2245) );
  OAI221_X1 U979 ( .B1(n17429), .B2(n18525), .C1(n17533), .C2(n18522), .A(
        n2248), .ZN(n2243) );
  NOR4_X1 U980 ( .A1(n2190), .A2(n2191), .A3(n2192), .A4(n2193), .ZN(n2189) );
  OAI221_X1 U981 ( .B1(n17750), .B2(n18513), .C1(n18261), .C2(n18510), .A(
        n2211), .ZN(n2190) );
  OAI221_X1 U982 ( .B1(n17366), .B2(n18548), .C1(n17621), .C2(n18545), .A(
        n2196), .ZN(n2193) );
  OAI221_X1 U983 ( .B1(n17430), .B2(n18525), .C1(n17534), .C2(n18522), .A(
        n2206), .ZN(n2191) );
  AND3_X1 U984 ( .A1(ADD_RD1[1]), .A2(n18352), .A3(ADD_RD1[2]), .ZN(n3914) );
  AND3_X1 U985 ( .A1(n17839), .A2(n4553), .A3(ADD_RD2[1]), .ZN(n4535) );
  AND3_X1 U986 ( .A1(n18352), .A2(n3925), .A3(ADD_RD1[2]), .ZN(n3907) );
  AND3_X1 U987 ( .A1(ADD_RD2[1]), .A2(n17839), .A3(ADD_RD2[2]), .ZN(n4538) );
  OAI22_X1 U988 ( .A1(n17679), .A2(n18403), .B1(n18000), .B2(n18400), .ZN(
        n4105) );
  OAI22_X1 U989 ( .A1(n17680), .A2(n18403), .B1(n18001), .B2(n18400), .ZN(
        n4087) );
  OAI22_X1 U990 ( .A1(n17681), .A2(n18403), .B1(n18002), .B2(n18400), .ZN(
        n4069) );
  OAI22_X1 U991 ( .A1(n17682), .A2(n18403), .B1(n18003), .B2(n18400), .ZN(
        n4051) );
  OAI22_X1 U992 ( .A1(n17683), .A2(n18403), .B1(n18004), .B2(n18400), .ZN(
        n4033) );
  OAI22_X1 U993 ( .A1(n17684), .A2(n18403), .B1(n18005), .B2(n18400), .ZN(
        n4015) );
  OAI22_X1 U994 ( .A1(n17685), .A2(n18403), .B1(n18006), .B2(n18400), .ZN(
        n3997) );
  OAI22_X1 U995 ( .A1(n17686), .A2(n18403), .B1(n18007), .B2(n18400), .ZN(
        n3962) );
  OAI22_X1 U996 ( .A1(n17872), .A2(n18501), .B1(n17661), .B2(n18498), .ZN(
        n2367) );
  OAI22_X1 U997 ( .A1(n17873), .A2(n18501), .B1(n17662), .B2(n18498), .ZN(
        n2348) );
  OAI22_X1 U998 ( .A1(n17874), .A2(n18501), .B1(n17663), .B2(n18498), .ZN(
        n2329) );
  OAI22_X1 U999 ( .A1(n17875), .A2(n18501), .B1(n17664), .B2(n18498), .ZN(
        n2310) );
  OAI22_X1 U1000 ( .A1(n17876), .A2(n18501), .B1(n17665), .B2(n18498), .ZN(
        n2291) );
  OAI22_X1 U1001 ( .A1(n17877), .A2(n18501), .B1(n17666), .B2(n18498), .ZN(
        n2272) );
  OAI22_X1 U1002 ( .A1(n17878), .A2(n18501), .B1(n17667), .B2(n18498), .ZN(
        n2253) );
  OAI22_X1 U1003 ( .A1(n17879), .A2(n18501), .B1(n17668), .B2(n18498), .ZN(
        n2217) );
  OAI22_X1 U1004 ( .A1(n17527), .A2(n18397), .B1(n17968), .B2(n18394), .ZN(
        n4104) );
  OAI22_X1 U1005 ( .A1(n17528), .A2(n18397), .B1(n17969), .B2(n18394), .ZN(
        n4086) );
  OAI22_X1 U1006 ( .A1(n17529), .A2(n18397), .B1(n17970), .B2(n18394), .ZN(
        n4068) );
  OAI22_X1 U1007 ( .A1(n17530), .A2(n18397), .B1(n17971), .B2(n18394), .ZN(
        n4050) );
  OAI22_X1 U1008 ( .A1(n17531), .A2(n18397), .B1(n17972), .B2(n18394), .ZN(
        n4032) );
  OAI22_X1 U1009 ( .A1(n17532), .A2(n18397), .B1(n17973), .B2(n18394), .ZN(
        n4014) );
  OAI22_X1 U1010 ( .A1(n17533), .A2(n18397), .B1(n17974), .B2(n18394), .ZN(
        n3996) );
  OAI22_X1 U1011 ( .A1(n17534), .A2(n18397), .B1(n17975), .B2(n18394), .ZN(
        n3961) );
  OAI22_X1 U1012 ( .A1(n17606), .A2(n18495), .B1(n17327), .B2(n18492), .ZN(
        n2366) );
  OAI22_X1 U1013 ( .A1(n17607), .A2(n18495), .B1(n17328), .B2(n18492), .ZN(
        n2347) );
  OAI22_X1 U1014 ( .A1(n17608), .A2(n18495), .B1(n17329), .B2(n18492), .ZN(
        n2328) );
  OAI22_X1 U1015 ( .A1(n17609), .A2(n18495), .B1(n17330), .B2(n18492), .ZN(
        n2309) );
  OAI22_X1 U1016 ( .A1(n17610), .A2(n18495), .B1(n17331), .B2(n18492), .ZN(
        n2290) );
  OAI22_X1 U1017 ( .A1(n17611), .A2(n18495), .B1(n17332), .B2(n18492), .ZN(
        n2271) );
  OAI22_X1 U1018 ( .A1(n17612), .A2(n18495), .B1(n17333), .B2(n18492), .ZN(
        n2252) );
  OAI22_X1 U1019 ( .A1(n17613), .A2(n18495), .B1(n17334), .B2(n18492), .ZN(
        n2216) );
  OAI22_X1 U1020 ( .A1(n17840), .A2(n18468), .B1(n17391), .B2(n18465), .ZN(
        n2368) );
  OAI22_X1 U1021 ( .A1(n17841), .A2(n18468), .B1(n17392), .B2(n18465), .ZN(
        n2349) );
  OAI22_X1 U1022 ( .A1(n17842), .A2(n18468), .B1(n17393), .B2(n18465), .ZN(
        n2330) );
  OAI22_X1 U1023 ( .A1(n17843), .A2(n18468), .B1(n17394), .B2(n18465), .ZN(
        n2311) );
  OAI22_X1 U1024 ( .A1(n17844), .A2(n18468), .B1(n17395), .B2(n18465), .ZN(
        n2292) );
  OAI22_X1 U1025 ( .A1(n17845), .A2(n18468), .B1(n17396), .B2(n18465), .ZN(
        n2273) );
  OAI22_X1 U1026 ( .A1(n17846), .A2(n18468), .B1(n17397), .B2(n18465), .ZN(
        n2254) );
  OAI22_X1 U1027 ( .A1(n17847), .A2(n18468), .B1(n17398), .B2(n18465), .ZN(
        n2229) );
  OAI22_X1 U1028 ( .A1(n17359), .A2(n18370), .B1(n18064), .B2(n18367), .ZN(
        n4106) );
  OAI22_X1 U1029 ( .A1(n17936), .A2(n18358), .B1(n17614), .B2(n18355), .ZN(
        n4107) );
  OAI22_X1 U1030 ( .A1(n17360), .A2(n18370), .B1(n18065), .B2(n18367), .ZN(
        n4088) );
  OAI22_X1 U1031 ( .A1(n17937), .A2(n18358), .B1(n17615), .B2(n18355), .ZN(
        n4089) );
  OAI22_X1 U1032 ( .A1(n17361), .A2(n18370), .B1(n18066), .B2(n18367), .ZN(
        n4070) );
  OAI22_X1 U1033 ( .A1(n17938), .A2(n18358), .B1(n17616), .B2(n18355), .ZN(
        n4071) );
  OAI22_X1 U1034 ( .A1(n17362), .A2(n18370), .B1(n18067), .B2(n18367), .ZN(
        n4052) );
  OAI22_X1 U1035 ( .A1(n17939), .A2(n18358), .B1(n17617), .B2(n18355), .ZN(
        n4053) );
  OAI22_X1 U1036 ( .A1(n17363), .A2(n18370), .B1(n18068), .B2(n18367), .ZN(
        n4034) );
  OAI22_X1 U1037 ( .A1(n17940), .A2(n18358), .B1(n17618), .B2(n18355), .ZN(
        n4035) );
  OAI22_X1 U1038 ( .A1(n17364), .A2(n18370), .B1(n18069), .B2(n18367), .ZN(
        n4016) );
  OAI22_X1 U1039 ( .A1(n17941), .A2(n18358), .B1(n17619), .B2(n18355), .ZN(
        n4017) );
  OAI22_X1 U1040 ( .A1(n17365), .A2(n18370), .B1(n18070), .B2(n18367), .ZN(
        n3998) );
  OAI22_X1 U1041 ( .A1(n17942), .A2(n18358), .B1(n17620), .B2(n18355), .ZN(
        n3999) );
  OAI22_X1 U1042 ( .A1(n17366), .A2(n18370), .B1(n18071), .B2(n18367), .ZN(
        n3974) );
  OAI22_X1 U1043 ( .A1(n17943), .A2(n18358), .B1(n17621), .B2(n18355), .ZN(
        n3979) );
  OAI22_X1 U1044 ( .A1(n17487), .A2(n18456), .B1(n18072), .B2(n18453), .ZN(
        n2369) );
  OAI22_X1 U1045 ( .A1(n17488), .A2(n18456), .B1(n18073), .B2(n18453), .ZN(
        n2350) );
  OAI22_X1 U1046 ( .A1(n17489), .A2(n18456), .B1(n18074), .B2(n18453), .ZN(
        n2331) );
  OAI22_X1 U1047 ( .A1(n17490), .A2(n18456), .B1(n18075), .B2(n18453), .ZN(
        n2312) );
  OAI22_X1 U1048 ( .A1(n17491), .A2(n18456), .B1(n18076), .B2(n18453), .ZN(
        n2293) );
  OAI22_X1 U1049 ( .A1(n17492), .A2(n18456), .B1(n18077), .B2(n18453), .ZN(
        n2274) );
  OAI22_X1 U1050 ( .A1(n17493), .A2(n18456), .B1(n18078), .B2(n18453), .ZN(
        n2255) );
  OAI22_X1 U1051 ( .A1(n17494), .A2(n18456), .B1(n18079), .B2(n18453), .ZN(
        n2234) );
  OAI22_X1 U1052 ( .A1(n17687), .A2(n18401), .B1(n18016), .B2(n18398), .ZN(
        n4549) );
  OAI22_X1 U1053 ( .A1(n17688), .A2(n18401), .B1(n18017), .B2(n18398), .ZN(
        n4519) );
  OAI22_X1 U1054 ( .A1(n17689), .A2(n18401), .B1(n18022), .B2(n18398), .ZN(
        n4501) );
  OAI22_X1 U1055 ( .A1(n17691), .A2(n18401), .B1(n18023), .B2(n18398), .ZN(
        n4483) );
  OAI22_X1 U1056 ( .A1(n17690), .A2(n18401), .B1(n18018), .B2(n18398), .ZN(
        n4465) );
  OAI22_X1 U1057 ( .A1(n17692), .A2(n18401), .B1(n18024), .B2(n18398), .ZN(
        n4447) );
  OAI22_X1 U1058 ( .A1(n17693), .A2(n18401), .B1(n18025), .B2(n18398), .ZN(
        n4429) );
  OAI22_X1 U1059 ( .A1(n17694), .A2(n18401), .B1(n18026), .B2(n18398), .ZN(
        n4411) );
  OAI22_X1 U1060 ( .A1(n17695), .A2(n18401), .B1(n18027), .B2(n18398), .ZN(
        n4393) );
  OAI22_X1 U1061 ( .A1(n17696), .A2(n18401), .B1(n18028), .B2(n18398), .ZN(
        n4375) );
  OAI22_X1 U1062 ( .A1(n17697), .A2(n18401), .B1(n18029), .B2(n18398), .ZN(
        n4357) );
  OAI22_X1 U1063 ( .A1(n17698), .A2(n18401), .B1(n18030), .B2(n18398), .ZN(
        n4339) );
  OAI22_X1 U1064 ( .A1(n17699), .A2(n18402), .B1(n18031), .B2(n18399), .ZN(
        n4321) );
  OAI22_X1 U1065 ( .A1(n17700), .A2(n18402), .B1(n18032), .B2(n18399), .ZN(
        n4303) );
  OAI22_X1 U1066 ( .A1(n17701), .A2(n18402), .B1(n18033), .B2(n18399), .ZN(
        n4285) );
  OAI22_X1 U1067 ( .A1(n17702), .A2(n18402), .B1(n18034), .B2(n18399), .ZN(
        n4267) );
  OAI22_X1 U1068 ( .A1(n17703), .A2(n18402), .B1(n18035), .B2(n18399), .ZN(
        n4249) );
  OAI22_X1 U1069 ( .A1(n17704), .A2(n18402), .B1(n18036), .B2(n18399), .ZN(
        n4231) );
  OAI22_X1 U1070 ( .A1(n17705), .A2(n18402), .B1(n18037), .B2(n18399), .ZN(
        n4213) );
  OAI22_X1 U1071 ( .A1(n17706), .A2(n18402), .B1(n18038), .B2(n18399), .ZN(
        n4195) );
  OAI22_X1 U1072 ( .A1(n17707), .A2(n18402), .B1(n18039), .B2(n18399), .ZN(
        n4177) );
  OAI22_X1 U1073 ( .A1(n17708), .A2(n18402), .B1(n18040), .B2(n18399), .ZN(
        n4159) );
  OAI22_X1 U1074 ( .A1(n17709), .A2(n18402), .B1(n18041), .B2(n18399), .ZN(
        n4141) );
  OAI22_X1 U1075 ( .A1(n17710), .A2(n18402), .B1(n18042), .B2(n18399), .ZN(
        n4123) );
  OAI22_X1 U1076 ( .A1(n17880), .A2(n18499), .B1(n17638), .B2(n18496), .ZN(
        n3923) );
  OAI22_X1 U1077 ( .A1(n17883), .A2(n18499), .B1(n17639), .B2(n18496), .ZN(
        n3892) );
  OAI22_X1 U1078 ( .A1(n17881), .A2(n18499), .B1(n17678), .B2(n18496), .ZN(
        n3873) );
  OAI22_X1 U1079 ( .A1(n17882), .A2(n18499), .B1(n17640), .B2(n18496), .ZN(
        n3854) );
  OAI22_X1 U1080 ( .A1(n17884), .A2(n18499), .B1(n17641), .B2(n18496), .ZN(
        n2747) );
  OAI22_X1 U1081 ( .A1(n17885), .A2(n18499), .B1(n17642), .B2(n18496), .ZN(
        n2728) );
  OAI22_X1 U1082 ( .A1(n17886), .A2(n18499), .B1(n17643), .B2(n18496), .ZN(
        n2709) );
  OAI22_X1 U1083 ( .A1(n17887), .A2(n18499), .B1(n17644), .B2(n18496), .ZN(
        n2690) );
  OAI22_X1 U1084 ( .A1(n17888), .A2(n18499), .B1(n17645), .B2(n18496), .ZN(
        n2671) );
  OAI22_X1 U1085 ( .A1(n17889), .A2(n18499), .B1(n17646), .B2(n18496), .ZN(
        n2652) );
  OAI22_X1 U1086 ( .A1(n17890), .A2(n18499), .B1(n17647), .B2(n18496), .ZN(
        n2633) );
  OAI22_X1 U1087 ( .A1(n17891), .A2(n18499), .B1(n17648), .B2(n18496), .ZN(
        n2614) );
  OAI22_X1 U1088 ( .A1(n17892), .A2(n18500), .B1(n17649), .B2(n18497), .ZN(
        n2595) );
  OAI22_X1 U1089 ( .A1(n17893), .A2(n18500), .B1(n17650), .B2(n18497), .ZN(
        n2576) );
  OAI22_X1 U1090 ( .A1(n17894), .A2(n18500), .B1(n17651), .B2(n18497), .ZN(
        n2557) );
  OAI22_X1 U1091 ( .A1(n17895), .A2(n18500), .B1(n17652), .B2(n18497), .ZN(
        n2538) );
  OAI22_X1 U1092 ( .A1(n17896), .A2(n18500), .B1(n17653), .B2(n18497), .ZN(
        n2519) );
  OAI22_X1 U1093 ( .A1(n17897), .A2(n18500), .B1(n17654), .B2(n18497), .ZN(
        n2500) );
  OAI22_X1 U1094 ( .A1(n17898), .A2(n18500), .B1(n17655), .B2(n18497), .ZN(
        n2481) );
  OAI22_X1 U1095 ( .A1(n17899), .A2(n18500), .B1(n17656), .B2(n18497), .ZN(
        n2462) );
  OAI22_X1 U1096 ( .A1(n17900), .A2(n18500), .B1(n17657), .B2(n18497), .ZN(
        n2443) );
  OAI22_X1 U1097 ( .A1(n17901), .A2(n18500), .B1(n17658), .B2(n18497), .ZN(
        n2424) );
  OAI22_X1 U1098 ( .A1(n17902), .A2(n18500), .B1(n17659), .B2(n18497), .ZN(
        n2405) );
  OAI22_X1 U1099 ( .A1(n17903), .A2(n18500), .B1(n17660), .B2(n18497), .ZN(
        n2386) );
  OAI22_X1 U1100 ( .A1(n17904), .A2(n18391), .B1(n17327), .B2(n18388), .ZN(
        n4103) );
  OAI22_X1 U1101 ( .A1(n17905), .A2(n18391), .B1(n17328), .B2(n18388), .ZN(
        n4085) );
  OAI22_X1 U1102 ( .A1(n17906), .A2(n18391), .B1(n17329), .B2(n18388), .ZN(
        n4067) );
  OAI22_X1 U1103 ( .A1(n17907), .A2(n18391), .B1(n17330), .B2(n18388), .ZN(
        n4049) );
  OAI22_X1 U1104 ( .A1(n17908), .A2(n18391), .B1(n17331), .B2(n18388), .ZN(
        n4031) );
  OAI22_X1 U1105 ( .A1(n17909), .A2(n18391), .B1(n17332), .B2(n18388), .ZN(
        n4013) );
  OAI22_X1 U1106 ( .A1(n17910), .A2(n18391), .B1(n17333), .B2(n18388), .ZN(
        n3995) );
  OAI22_X1 U1107 ( .A1(n17911), .A2(n18391), .B1(n17334), .B2(n18388), .ZN(
        n3960) );
  OAI22_X1 U1108 ( .A1(n17519), .A2(n18489), .B1(n18008), .B2(n18486), .ZN(
        n2365) );
  OAI22_X1 U1109 ( .A1(n17520), .A2(n18489), .B1(n18009), .B2(n18486), .ZN(
        n2346) );
  OAI22_X1 U1110 ( .A1(n17521), .A2(n18489), .B1(n18010), .B2(n18486), .ZN(
        n2327) );
  OAI22_X1 U1111 ( .A1(n17522), .A2(n18489), .B1(n18011), .B2(n18486), .ZN(
        n2308) );
  OAI22_X1 U1112 ( .A1(n17523), .A2(n18489), .B1(n18012), .B2(n18486), .ZN(
        n2289) );
  OAI22_X1 U1113 ( .A1(n17524), .A2(n18489), .B1(n18013), .B2(n18486), .ZN(
        n2270) );
  OAI22_X1 U1114 ( .A1(n17525), .A2(n18489), .B1(n18014), .B2(n18486), .ZN(
        n2251) );
  OAI22_X1 U1115 ( .A1(n17526), .A2(n18489), .B1(n18015), .B2(n18486), .ZN(
        n2215) );
  OAI22_X1 U1116 ( .A1(n17537), .A2(n18395), .B1(n17979), .B2(n18392), .ZN(
        n4548) );
  OAI22_X1 U1117 ( .A1(n17562), .A2(n18395), .B1(n17980), .B2(n18392), .ZN(
        n4518) );
  OAI22_X1 U1118 ( .A1(n17538), .A2(n18395), .B1(n17976), .B2(n18392), .ZN(
        n4500) );
  OAI22_X1 U1119 ( .A1(n17563), .A2(n18395), .B1(n17977), .B2(n18392), .ZN(
        n4482) );
  OAI22_X1 U1120 ( .A1(n17539), .A2(n18395), .B1(n17978), .B2(n18392), .ZN(
        n4464) );
  OAI22_X1 U1121 ( .A1(n17564), .A2(n18395), .B1(n17981), .B2(n18392), .ZN(
        n4446) );
  OAI22_X1 U1122 ( .A1(n17565), .A2(n18395), .B1(n17982), .B2(n18392), .ZN(
        n4428) );
  OAI22_X1 U1123 ( .A1(n17566), .A2(n18395), .B1(n17983), .B2(n18392), .ZN(
        n4410) );
  OAI22_X1 U1124 ( .A1(n17567), .A2(n18395), .B1(n17984), .B2(n18392), .ZN(
        n4392) );
  OAI22_X1 U1125 ( .A1(n17568), .A2(n18395), .B1(n17985), .B2(n18392), .ZN(
        n4374) );
  OAI22_X1 U1126 ( .A1(n17569), .A2(n18395), .B1(n17986), .B2(n18392), .ZN(
        n4356) );
  OAI22_X1 U1127 ( .A1(n17570), .A2(n18395), .B1(n17987), .B2(n18392), .ZN(
        n4338) );
  OAI22_X1 U1128 ( .A1(n17571), .A2(n18396), .B1(n17988), .B2(n18393), .ZN(
        n4320) );
  OAI22_X1 U1129 ( .A1(n17572), .A2(n18396), .B1(n17989), .B2(n18393), .ZN(
        n4302) );
  OAI22_X1 U1130 ( .A1(n17573), .A2(n18396), .B1(n17990), .B2(n18393), .ZN(
        n4284) );
  OAI22_X1 U1131 ( .A1(n17574), .A2(n18396), .B1(n17991), .B2(n18393), .ZN(
        n4266) );
  OAI22_X1 U1132 ( .A1(n17575), .A2(n18396), .B1(n17992), .B2(n18393), .ZN(
        n4248) );
  OAI22_X1 U1133 ( .A1(n17576), .A2(n18396), .B1(n17993), .B2(n18393), .ZN(
        n4230) );
  OAI22_X1 U1134 ( .A1(n17577), .A2(n18396), .B1(n17994), .B2(n18393), .ZN(
        n4212) );
  OAI22_X1 U1135 ( .A1(n17578), .A2(n18396), .B1(n17995), .B2(n18393), .ZN(
        n4194) );
  OAI22_X1 U1136 ( .A1(n17579), .A2(n18396), .B1(n17996), .B2(n18393), .ZN(
        n4176) );
  OAI22_X1 U1137 ( .A1(n17580), .A2(n18396), .B1(n17997), .B2(n18393), .ZN(
        n4158) );
  OAI22_X1 U1138 ( .A1(n17581), .A2(n18396), .B1(n17998), .B2(n18393), .ZN(
        n4140) );
  OAI22_X1 U1139 ( .A1(n17582), .A2(n18396), .B1(n17999), .B2(n18393), .ZN(
        n4122) );
  OAI22_X1 U1140 ( .A1(n17583), .A2(n18493), .B1(n17335), .B2(n18490), .ZN(
        n3922) );
  OAI22_X1 U1141 ( .A1(n17677), .A2(n18493), .B1(n17338), .B2(n18490), .ZN(
        n3891) );
  OAI22_X1 U1142 ( .A1(n17584), .A2(n18493), .B1(n17339), .B2(n18490), .ZN(
        n3872) );
  OAI22_X1 U1143 ( .A1(n17585), .A2(n18493), .B1(n17336), .B2(n18490), .ZN(
        n3853) );
  OAI22_X1 U1144 ( .A1(n17586), .A2(n18493), .B1(n17337), .B2(n18490), .ZN(
        n2746) );
  OAI22_X1 U1145 ( .A1(n17587), .A2(n18493), .B1(n17340), .B2(n18490), .ZN(
        n2727) );
  OAI22_X1 U1146 ( .A1(n17588), .A2(n18493), .B1(n17341), .B2(n18490), .ZN(
        n2708) );
  OAI22_X1 U1147 ( .A1(n17589), .A2(n18493), .B1(n17342), .B2(n18490), .ZN(
        n2689) );
  OAI22_X1 U1148 ( .A1(n17590), .A2(n18493), .B1(n17343), .B2(n18490), .ZN(
        n2670) );
  OAI22_X1 U1149 ( .A1(n17591), .A2(n18493), .B1(n17344), .B2(n18490), .ZN(
        n2651) );
  OAI22_X1 U1150 ( .A1(n17592), .A2(n18493), .B1(n17345), .B2(n18490), .ZN(
        n2632) );
  OAI22_X1 U1151 ( .A1(n17593), .A2(n18493), .B1(n17346), .B2(n18490), .ZN(
        n2613) );
  OAI22_X1 U1152 ( .A1(n17594), .A2(n18494), .B1(n17347), .B2(n18491), .ZN(
        n2594) );
  OAI22_X1 U1153 ( .A1(n17595), .A2(n18494), .B1(n17348), .B2(n18491), .ZN(
        n2575) );
  OAI22_X1 U1154 ( .A1(n17596), .A2(n18494), .B1(n17349), .B2(n18491), .ZN(
        n2556) );
  OAI22_X1 U1155 ( .A1(n17597), .A2(n18494), .B1(n17350), .B2(n18491), .ZN(
        n2537) );
  OAI22_X1 U1156 ( .A1(n17598), .A2(n18494), .B1(n17351), .B2(n18491), .ZN(
        n2518) );
  OAI22_X1 U1157 ( .A1(n17599), .A2(n18494), .B1(n17352), .B2(n18491), .ZN(
        n2499) );
  OAI22_X1 U1158 ( .A1(n17600), .A2(n18494), .B1(n17353), .B2(n18491), .ZN(
        n2480) );
  OAI22_X1 U1159 ( .A1(n17601), .A2(n18494), .B1(n17354), .B2(n18491), .ZN(
        n2461) );
  OAI22_X1 U1160 ( .A1(n17602), .A2(n18494), .B1(n17355), .B2(n18491), .ZN(
        n2442) );
  OAI22_X1 U1161 ( .A1(n17603), .A2(n18494), .B1(n17356), .B2(n18491), .ZN(
        n2423) );
  OAI22_X1 U1162 ( .A1(n17604), .A2(n18494), .B1(n17357), .B2(n18491), .ZN(
        n2404) );
  OAI22_X1 U1163 ( .A1(n17605), .A2(n18494), .B1(n17358), .B2(n18491), .ZN(
        n2385) );
  OAI22_X1 U1164 ( .A1(n17383), .A2(n18368), .B1(n18080), .B2(n18365), .ZN(
        n4554) );
  OAI22_X1 U1165 ( .A1(n17944), .A2(n18356), .B1(n17669), .B2(n18353), .ZN(
        n4555) );
  OAI22_X1 U1166 ( .A1(n17384), .A2(n18368), .B1(n18081), .B2(n18365), .ZN(
        n4520) );
  OAI22_X1 U1167 ( .A1(n17945), .A2(n18356), .B1(n17670), .B2(n18353), .ZN(
        n4521) );
  OAI22_X1 U1168 ( .A1(n17385), .A2(n18368), .B1(n18082), .B2(n18365), .ZN(
        n4502) );
  OAI22_X1 U1169 ( .A1(n17946), .A2(n18356), .B1(n17671), .B2(n18353), .ZN(
        n4503) );
  OAI22_X1 U1170 ( .A1(n17386), .A2(n18368), .B1(n18083), .B2(n18365), .ZN(
        n4484) );
  OAI22_X1 U1171 ( .A1(n17947), .A2(n18356), .B1(n17672), .B2(n18353), .ZN(
        n4485) );
  OAI22_X1 U1172 ( .A1(n17387), .A2(n18368), .B1(n18086), .B2(n18365), .ZN(
        n4466) );
  OAI22_X1 U1173 ( .A1(n17948), .A2(n18356), .B1(n17673), .B2(n18353), .ZN(
        n4467) );
  OAI22_X1 U1174 ( .A1(n17388), .A2(n18368), .B1(n18087), .B2(n18365), .ZN(
        n4448) );
  OAI22_X1 U1175 ( .A1(n17949), .A2(n18356), .B1(n17674), .B2(n18353), .ZN(
        n4449) );
  OAI22_X1 U1176 ( .A1(n17389), .A2(n18368), .B1(n18088), .B2(n18365), .ZN(
        n4430) );
  OAI22_X1 U1177 ( .A1(n17950), .A2(n18356), .B1(n17675), .B2(n18353), .ZN(
        n4431) );
  OAI22_X1 U1178 ( .A1(n17390), .A2(n18368), .B1(n18089), .B2(n18365), .ZN(
        n4412) );
  OAI22_X1 U1179 ( .A1(n17951), .A2(n18356), .B1(n17676), .B2(n18353), .ZN(
        n4413) );
  OAI22_X1 U1180 ( .A1(n17367), .A2(n18368), .B1(n18090), .B2(n18365), .ZN(
        n4394) );
  OAI22_X1 U1181 ( .A1(n17952), .A2(n18356), .B1(n17622), .B2(n18353), .ZN(
        n4395) );
  OAI22_X1 U1182 ( .A1(n17368), .A2(n18368), .B1(n18091), .B2(n18365), .ZN(
        n4376) );
  OAI22_X1 U1183 ( .A1(n17953), .A2(n18356), .B1(n17623), .B2(n18353), .ZN(
        n4377) );
  OAI22_X1 U1184 ( .A1(n17369), .A2(n18368), .B1(n18092), .B2(n18365), .ZN(
        n4358) );
  OAI22_X1 U1185 ( .A1(n17954), .A2(n18356), .B1(n17624), .B2(n18353), .ZN(
        n4359) );
  OAI22_X1 U1186 ( .A1(n17370), .A2(n18368), .B1(n18093), .B2(n18365), .ZN(
        n4340) );
  OAI22_X1 U1187 ( .A1(n17955), .A2(n18356), .B1(n17625), .B2(n18353), .ZN(
        n4341) );
  OAI22_X1 U1188 ( .A1(n17371), .A2(n18369), .B1(n18094), .B2(n18366), .ZN(
        n4322) );
  OAI22_X1 U1189 ( .A1(n17956), .A2(n18357), .B1(n17626), .B2(n18354), .ZN(
        n4323) );
  OAI22_X1 U1190 ( .A1(n17372), .A2(n18369), .B1(n18095), .B2(n18366), .ZN(
        n4304) );
  OAI22_X1 U1191 ( .A1(n17957), .A2(n18357), .B1(n17627), .B2(n18354), .ZN(
        n4305) );
  OAI22_X1 U1192 ( .A1(n17373), .A2(n18369), .B1(n18096), .B2(n18366), .ZN(
        n4286) );
  OAI22_X1 U1193 ( .A1(n17958), .A2(n18357), .B1(n17628), .B2(n18354), .ZN(
        n4287) );
  OAI22_X1 U1194 ( .A1(n17374), .A2(n18369), .B1(n18097), .B2(n18366), .ZN(
        n4268) );
  OAI22_X1 U1195 ( .A1(n17959), .A2(n18357), .B1(n17629), .B2(n18354), .ZN(
        n4269) );
  OAI22_X1 U1196 ( .A1(n17375), .A2(n18369), .B1(n18098), .B2(n18366), .ZN(
        n4250) );
  OAI22_X1 U1197 ( .A1(n17960), .A2(n18357), .B1(n17630), .B2(n18354), .ZN(
        n4251) );
  OAI22_X1 U1198 ( .A1(n17376), .A2(n18369), .B1(n18099), .B2(n18366), .ZN(
        n4232) );
  OAI22_X1 U1199 ( .A1(n17961), .A2(n18357), .B1(n17631), .B2(n18354), .ZN(
        n4233) );
  OAI22_X1 U1200 ( .A1(n17377), .A2(n18369), .B1(n18100), .B2(n18366), .ZN(
        n4214) );
  OAI22_X1 U1201 ( .A1(n17962), .A2(n18357), .B1(n17632), .B2(n18354), .ZN(
        n4215) );
  OAI22_X1 U1202 ( .A1(n17378), .A2(n18369), .B1(n18101), .B2(n18366), .ZN(
        n4196) );
  OAI22_X1 U1203 ( .A1(n17963), .A2(n18357), .B1(n17633), .B2(n18354), .ZN(
        n4197) );
  OAI22_X1 U1204 ( .A1(n17379), .A2(n18369), .B1(n18102), .B2(n18366), .ZN(
        n4178) );
  OAI22_X1 U1205 ( .A1(n17964), .A2(n18357), .B1(n17634), .B2(n18354), .ZN(
        n4179) );
  OAI22_X1 U1206 ( .A1(n17380), .A2(n18369), .B1(n18103), .B2(n18366), .ZN(
        n4160) );
  OAI22_X1 U1207 ( .A1(n17965), .A2(n18357), .B1(n17635), .B2(n18354), .ZN(
        n4161) );
  OAI22_X1 U1208 ( .A1(n17381), .A2(n18369), .B1(n18104), .B2(n18366), .ZN(
        n4142) );
  OAI22_X1 U1209 ( .A1(n17966), .A2(n18357), .B1(n17636), .B2(n18354), .ZN(
        n4143) );
  OAI22_X1 U1210 ( .A1(n17382), .A2(n18369), .B1(n18105), .B2(n18366), .ZN(
        n4124) );
  OAI22_X1 U1211 ( .A1(n17967), .A2(n18357), .B1(n17637), .B2(n18354), .ZN(
        n4125) );
  OAI22_X1 U1212 ( .A1(n17518), .A2(n18454), .B1(n18106), .B2(n18451), .ZN(
        n3930) );
  OAI22_X1 U1213 ( .A1(n17848), .A2(n18466), .B1(n17402), .B2(n18463), .ZN(
        n3927) );
  OAI22_X1 U1214 ( .A1(n17495), .A2(n18454), .B1(n18107), .B2(n18451), .ZN(
        n3894) );
  OAI22_X1 U1215 ( .A1(n17849), .A2(n18466), .B1(n17399), .B2(n18463), .ZN(
        n3893) );
  OAI22_X1 U1216 ( .A1(n17496), .A2(n18454), .B1(n18084), .B2(n18451), .ZN(
        n3875) );
  OAI22_X1 U1217 ( .A1(n17850), .A2(n18466), .B1(n17400), .B2(n18463), .ZN(
        n3874) );
  OAI22_X1 U1218 ( .A1(n17497), .A2(n18454), .B1(n18108), .B2(n18451), .ZN(
        n3856) );
  OAI22_X1 U1219 ( .A1(n17851), .A2(n18466), .B1(n17403), .B2(n18463), .ZN(
        n3855) );
  OAI22_X1 U1220 ( .A1(n17498), .A2(n18454), .B1(n18085), .B2(n18451), .ZN(
        n2749) );
  OAI22_X1 U1221 ( .A1(n17852), .A2(n18466), .B1(n17401), .B2(n18463), .ZN(
        n2748) );
  OAI22_X1 U1222 ( .A1(n17499), .A2(n18454), .B1(n18109), .B2(n18451), .ZN(
        n2730) );
  OAI22_X1 U1223 ( .A1(n17853), .A2(n18466), .B1(n17404), .B2(n18463), .ZN(
        n2729) );
  OAI22_X1 U1224 ( .A1(n17500), .A2(n18454), .B1(n18110), .B2(n18451), .ZN(
        n2711) );
  OAI22_X1 U1225 ( .A1(n17854), .A2(n18466), .B1(n17405), .B2(n18463), .ZN(
        n2710) );
  OAI22_X1 U1226 ( .A1(n17501), .A2(n18454), .B1(n18111), .B2(n18451), .ZN(
        n2692) );
  OAI22_X1 U1227 ( .A1(n17855), .A2(n18466), .B1(n17406), .B2(n18463), .ZN(
        n2691) );
  OAI22_X1 U1228 ( .A1(n17502), .A2(n18454), .B1(n18112), .B2(n18451), .ZN(
        n2673) );
  OAI22_X1 U1229 ( .A1(n17856), .A2(n18466), .B1(n17407), .B2(n18463), .ZN(
        n2672) );
  OAI22_X1 U1230 ( .A1(n17503), .A2(n18454), .B1(n18113), .B2(n18451), .ZN(
        n2654) );
  OAI22_X1 U1231 ( .A1(n17857), .A2(n18466), .B1(n17408), .B2(n18463), .ZN(
        n2653) );
  OAI22_X1 U1232 ( .A1(n17504), .A2(n18454), .B1(n18114), .B2(n18451), .ZN(
        n2635) );
  OAI22_X1 U1233 ( .A1(n17858), .A2(n18466), .B1(n17409), .B2(n18463), .ZN(
        n2634) );
  OAI22_X1 U1234 ( .A1(n17505), .A2(n18454), .B1(n18115), .B2(n18451), .ZN(
        n2616) );
  OAI22_X1 U1235 ( .A1(n17859), .A2(n18466), .B1(n17410), .B2(n18463), .ZN(
        n2615) );
  OAI22_X1 U1236 ( .A1(n17506), .A2(n18455), .B1(n18116), .B2(n18452), .ZN(
        n2597) );
  OAI22_X1 U1237 ( .A1(n17860), .A2(n18467), .B1(n17411), .B2(n18464), .ZN(
        n2596) );
  OAI22_X1 U1238 ( .A1(n17507), .A2(n18455), .B1(n18117), .B2(n18452), .ZN(
        n2578) );
  OAI22_X1 U1239 ( .A1(n17861), .A2(n18467), .B1(n17412), .B2(n18464), .ZN(
        n2577) );
  OAI22_X1 U1240 ( .A1(n17508), .A2(n18455), .B1(n18118), .B2(n18452), .ZN(
        n2559) );
  OAI22_X1 U1241 ( .A1(n17862), .A2(n18467), .B1(n17413), .B2(n18464), .ZN(
        n2558) );
  OAI22_X1 U1242 ( .A1(n17509), .A2(n18455), .B1(n18119), .B2(n18452), .ZN(
        n2540) );
  OAI22_X1 U1243 ( .A1(n17863), .A2(n18467), .B1(n17414), .B2(n18464), .ZN(
        n2539) );
  OAI22_X1 U1244 ( .A1(n17510), .A2(n18455), .B1(n18120), .B2(n18452), .ZN(
        n2521) );
  OAI22_X1 U1245 ( .A1(n17864), .A2(n18467), .B1(n17415), .B2(n18464), .ZN(
        n2520) );
  OAI22_X1 U1246 ( .A1(n17511), .A2(n18455), .B1(n18121), .B2(n18452), .ZN(
        n2502) );
  OAI22_X1 U1247 ( .A1(n17865), .A2(n18467), .B1(n17416), .B2(n18464), .ZN(
        n2501) );
  OAI22_X1 U1248 ( .A1(n17512), .A2(n18455), .B1(n18122), .B2(n18452), .ZN(
        n2483) );
  OAI22_X1 U1249 ( .A1(n17866), .A2(n18467), .B1(n17417), .B2(n18464), .ZN(
        n2482) );
  OAI22_X1 U1250 ( .A1(n17513), .A2(n18455), .B1(n18123), .B2(n18452), .ZN(
        n2464) );
  OAI22_X1 U1251 ( .A1(n17867), .A2(n18467), .B1(n17418), .B2(n18464), .ZN(
        n2463) );
  OAI22_X1 U1252 ( .A1(n17514), .A2(n18455), .B1(n18124), .B2(n18452), .ZN(
        n2445) );
  OAI22_X1 U1253 ( .A1(n17868), .A2(n18467), .B1(n17419), .B2(n18464), .ZN(
        n2444) );
  OAI22_X1 U1254 ( .A1(n17515), .A2(n18455), .B1(n18125), .B2(n18452), .ZN(
        n2426) );
  OAI22_X1 U1255 ( .A1(n17869), .A2(n18467), .B1(n17420), .B2(n18464), .ZN(
        n2425) );
  OAI22_X1 U1256 ( .A1(n17516), .A2(n18455), .B1(n18126), .B2(n18452), .ZN(
        n2407) );
  OAI22_X1 U1257 ( .A1(n17870), .A2(n18467), .B1(n17421), .B2(n18464), .ZN(
        n2406) );
  OAI22_X1 U1258 ( .A1(n17517), .A2(n18455), .B1(n18127), .B2(n18452), .ZN(
        n2388) );
  OAI22_X1 U1259 ( .A1(n17871), .A2(n18467), .B1(n17422), .B2(n18464), .ZN(
        n2387) );
  OAI22_X1 U1260 ( .A1(n17914), .A2(n18389), .B1(n17335), .B2(n18386), .ZN(
        n4547) );
  OAI22_X1 U1261 ( .A1(n17912), .A2(n18389), .B1(n17338), .B2(n18386), .ZN(
        n4517) );
  OAI22_X1 U1262 ( .A1(n17913), .A2(n18389), .B1(n17339), .B2(n18386), .ZN(
        n4499) );
  OAI22_X1 U1263 ( .A1(n17915), .A2(n18389), .B1(n17336), .B2(n18386), .ZN(
        n4481) );
  OAI22_X1 U1264 ( .A1(n17916), .A2(n18389), .B1(n17337), .B2(n18386), .ZN(
        n4463) );
  OAI22_X1 U1265 ( .A1(n17917), .A2(n18389), .B1(n17340), .B2(n18386), .ZN(
        n4445) );
  OAI22_X1 U1266 ( .A1(n17918), .A2(n18389), .B1(n17341), .B2(n18386), .ZN(
        n4427) );
  OAI22_X1 U1267 ( .A1(n17919), .A2(n18389), .B1(n17342), .B2(n18386), .ZN(
        n4409) );
  OAI22_X1 U1268 ( .A1(n17920), .A2(n18389), .B1(n17343), .B2(n18386), .ZN(
        n4391) );
  OAI22_X1 U1269 ( .A1(n17921), .A2(n18389), .B1(n17344), .B2(n18386), .ZN(
        n4373) );
  OAI22_X1 U1270 ( .A1(n17922), .A2(n18389), .B1(n17345), .B2(n18386), .ZN(
        n4355) );
  OAI22_X1 U1271 ( .A1(n17923), .A2(n18389), .B1(n17346), .B2(n18386), .ZN(
        n4337) );
  OAI22_X1 U1272 ( .A1(n17924), .A2(n18390), .B1(n17347), .B2(n18387), .ZN(
        n4319) );
  OAI22_X1 U1273 ( .A1(n17925), .A2(n18390), .B1(n17348), .B2(n18387), .ZN(
        n4301) );
  OAI22_X1 U1274 ( .A1(n17926), .A2(n18390), .B1(n17349), .B2(n18387), .ZN(
        n4283) );
  OAI22_X1 U1275 ( .A1(n17927), .A2(n18390), .B1(n17350), .B2(n18387), .ZN(
        n4265) );
  OAI22_X1 U1276 ( .A1(n17928), .A2(n18390), .B1(n17351), .B2(n18387), .ZN(
        n4247) );
  OAI22_X1 U1277 ( .A1(n17929), .A2(n18390), .B1(n17352), .B2(n18387), .ZN(
        n4229) );
  OAI22_X1 U1278 ( .A1(n17930), .A2(n18390), .B1(n17353), .B2(n18387), .ZN(
        n4211) );
  OAI22_X1 U1279 ( .A1(n17931), .A2(n18390), .B1(n17354), .B2(n18387), .ZN(
        n4193) );
  OAI22_X1 U1280 ( .A1(n17932), .A2(n18390), .B1(n17355), .B2(n18387), .ZN(
        n4175) );
  OAI22_X1 U1281 ( .A1(n17933), .A2(n18390), .B1(n17356), .B2(n18387), .ZN(
        n4157) );
  OAI22_X1 U1282 ( .A1(n17934), .A2(n18390), .B1(n17357), .B2(n18387), .ZN(
        n4139) );
  OAI22_X1 U1283 ( .A1(n17935), .A2(n18390), .B1(n17358), .B2(n18387), .ZN(
        n4121) );
  OAI22_X1 U1284 ( .A1(n17535), .A2(n18487), .B1(n18043), .B2(n18484), .ZN(
        n3921) );
  OAI22_X1 U1285 ( .A1(n17536), .A2(n18487), .B1(n18019), .B2(n18484), .ZN(
        n3890) );
  OAI22_X1 U1286 ( .A1(n17540), .A2(n18487), .B1(n18044), .B2(n18484), .ZN(
        n3871) );
  OAI22_X1 U1287 ( .A1(n17541), .A2(n18487), .B1(n18020), .B2(n18484), .ZN(
        n3852) );
  OAI22_X1 U1288 ( .A1(n17542), .A2(n18487), .B1(n18021), .B2(n18484), .ZN(
        n2745) );
  OAI22_X1 U1289 ( .A1(n17543), .A2(n18487), .B1(n18045), .B2(n18484), .ZN(
        n2726) );
  OAI22_X1 U1290 ( .A1(n17544), .A2(n18487), .B1(n18046), .B2(n18484), .ZN(
        n2707) );
  OAI22_X1 U1291 ( .A1(n17545), .A2(n18487), .B1(n18047), .B2(n18484), .ZN(
        n2688) );
  OAI22_X1 U1292 ( .A1(n17546), .A2(n18487), .B1(n18048), .B2(n18484), .ZN(
        n2669) );
  OAI22_X1 U1293 ( .A1(n17547), .A2(n18487), .B1(n18049), .B2(n18484), .ZN(
        n2650) );
  OAI22_X1 U1294 ( .A1(n17548), .A2(n18487), .B1(n18050), .B2(n18484), .ZN(
        n2631) );
  OAI22_X1 U1295 ( .A1(n17549), .A2(n18487), .B1(n18051), .B2(n18484), .ZN(
        n2612) );
  OAI22_X1 U1296 ( .A1(n17550), .A2(n18488), .B1(n18052), .B2(n18485), .ZN(
        n2593) );
  OAI22_X1 U1297 ( .A1(n17551), .A2(n18488), .B1(n18053), .B2(n18485), .ZN(
        n2574) );
  OAI22_X1 U1298 ( .A1(n17552), .A2(n18488), .B1(n18054), .B2(n18485), .ZN(
        n2555) );
  OAI22_X1 U1299 ( .A1(n17553), .A2(n18488), .B1(n18055), .B2(n18485), .ZN(
        n2536) );
  OAI22_X1 U1300 ( .A1(n17554), .A2(n18488), .B1(n18056), .B2(n18485), .ZN(
        n2517) );
  OAI22_X1 U1301 ( .A1(n17555), .A2(n18488), .B1(n18057), .B2(n18485), .ZN(
        n2498) );
  OAI22_X1 U1302 ( .A1(n17556), .A2(n18488), .B1(n18058), .B2(n18485), .ZN(
        n2479) );
  OAI22_X1 U1303 ( .A1(n17557), .A2(n18488), .B1(n18059), .B2(n18485), .ZN(
        n2460) );
  OAI22_X1 U1304 ( .A1(n17558), .A2(n18488), .B1(n18060), .B2(n18485), .ZN(
        n2441) );
  OAI22_X1 U1305 ( .A1(n17559), .A2(n18488), .B1(n18061), .B2(n18485), .ZN(
        n2422) );
  OAI22_X1 U1306 ( .A1(n17560), .A2(n18488), .B1(n18062), .B2(n18485), .ZN(
        n2403) );
  OAI22_X1 U1307 ( .A1(n17561), .A2(n18488), .B1(n18063), .B2(n18485), .ZN(
        n2384) );
  INV_X1 U1308 ( .A(ADD_RD1[3]), .ZN(n3928) );
  INV_X1 U1309 ( .A(ADD_RD1[0]), .ZN(n3929) );
  INV_X1 U1310 ( .A(ADD_RD1[4]), .ZN(n3926) );
  INV_X1 U1311 ( .A(ADD_RD1[1]), .ZN(n3925) );
  OAI21_X1 U1312 ( .B1(n1247), .B2(n2112), .A(n18997), .ZN(n2183) );
  OAI22_X1 U1313 ( .A1(n18570), .A2(n17518), .B1(n18561), .B2(n1136), .ZN(
        n2856) );
  OAI22_X1 U1314 ( .A1(n18584), .A2(n17677), .B1(n18575), .B2(n1134), .ZN(
        n2889) );
  OAI22_X1 U1315 ( .A1(n18610), .A2(n17678), .B1(n18601), .B2(n1132), .ZN(
        n2954) );
  OAI22_X1 U1316 ( .A1(n18657), .A2(n18286), .B1(n18648), .B2(n1130), .ZN(
        n3083) );
  OAI22_X1 U1317 ( .A1(n18748), .A2(n18287), .B1(n18739), .B2(n1128), .ZN(
        n3340) );
  BUF_X1 U1318 ( .A(n1126), .Z(n18905) );
  BUF_X1 U1319 ( .A(n1124), .Z(n18908) );
  BUF_X1 U1320 ( .A(n1122), .Z(n18911) );
  BUF_X1 U1321 ( .A(n1120), .Z(n18914) );
  BUF_X1 U1322 ( .A(n1118), .Z(n18917) );
  BUF_X1 U1323 ( .A(n1116), .Z(n18920) );
  BUF_X1 U1324 ( .A(n1114), .Z(n18923) );
  BUF_X1 U1325 ( .A(n1112), .Z(n18926) );
  BUF_X1 U1326 ( .A(n1110), .Z(n18929) );
  BUF_X1 U1327 ( .A(n1108), .Z(n18932) );
  BUF_X1 U1328 ( .A(n1106), .Z(n18935) );
  BUF_X1 U1329 ( .A(n1104), .Z(n18938) );
  BUF_X1 U1330 ( .A(n1102), .Z(n18941) );
  BUF_X1 U1331 ( .A(n1100), .Z(n18944) );
  BUF_X1 U1332 ( .A(n1098), .Z(n18947) );
  BUF_X1 U1333 ( .A(n1096), .Z(n18950) );
  BUF_X1 U1334 ( .A(n1094), .Z(n18953) );
  BUF_X1 U1335 ( .A(n1092), .Z(n18956) );
  BUF_X1 U1336 ( .A(n1090), .Z(n18959) );
  BUF_X1 U1337 ( .A(n1088), .Z(n18962) );
  BUF_X1 U1338 ( .A(n1086), .Z(n18965) );
  BUF_X1 U1339 ( .A(n1084), .Z(n18968) );
  BUF_X1 U1340 ( .A(n1082), .Z(n18971) );
  BUF_X1 U1341 ( .A(n1080), .Z(n18974) );
  BUF_X1 U1342 ( .A(n1126), .Z(n18904) );
  BUF_X1 U1343 ( .A(n1124), .Z(n18907) );
  BUF_X1 U1344 ( .A(n1122), .Z(n18910) );
  BUF_X1 U1345 ( .A(n1120), .Z(n18913) );
  BUF_X1 U1346 ( .A(n1118), .Z(n18916) );
  BUF_X1 U1347 ( .A(n1116), .Z(n18919) );
  BUF_X1 U1348 ( .A(n1114), .Z(n18922) );
  BUF_X1 U1349 ( .A(n1112), .Z(n18925) );
  BUF_X1 U1350 ( .A(n1110), .Z(n18928) );
  BUF_X1 U1351 ( .A(n1108), .Z(n18931) );
  BUF_X1 U1352 ( .A(n1106), .Z(n18934) );
  BUF_X1 U1353 ( .A(n1104), .Z(n18937) );
  BUF_X1 U1354 ( .A(n1102), .Z(n18940) );
  BUF_X1 U1355 ( .A(n1100), .Z(n18943) );
  BUF_X1 U1356 ( .A(n1098), .Z(n18946) );
  BUF_X1 U1357 ( .A(n1096), .Z(n18949) );
  BUF_X1 U1358 ( .A(n1094), .Z(n18952) );
  BUF_X1 U1359 ( .A(n1092), .Z(n18955) );
  BUF_X1 U1360 ( .A(n1090), .Z(n18958) );
  BUF_X1 U1361 ( .A(n1088), .Z(n18961) );
  BUF_X1 U1362 ( .A(n1086), .Z(n18964) );
  BUF_X1 U1363 ( .A(n1084), .Z(n18967) );
  BUF_X1 U1364 ( .A(n1082), .Z(n18970) );
  BUF_X1 U1365 ( .A(n1080), .Z(n18973) );
  BUF_X1 U1366 ( .A(n1078), .Z(n18977) );
  BUF_X1 U1367 ( .A(n1076), .Z(n18980) );
  BUF_X1 U1368 ( .A(n1073), .Z(n18992) );
  BUF_X1 U1369 ( .A(n1078), .Z(n18976) );
  BUF_X1 U1370 ( .A(n1076), .Z(n18979) );
  BUF_X1 U1371 ( .A(n1073), .Z(n18991) );
  BUF_X1 U1372 ( .A(RESET), .Z(n18995) );
  BUF_X1 U1373 ( .A(RESET), .Z(n18994) );
  BUF_X1 U1374 ( .A(n1126), .Z(n18906) );
  BUF_X1 U1375 ( .A(n1124), .Z(n18909) );
  BUF_X1 U1376 ( .A(n1122), .Z(n18912) );
  BUF_X1 U1377 ( .A(n1120), .Z(n18915) );
  BUF_X1 U1378 ( .A(n1118), .Z(n18918) );
  BUF_X1 U1379 ( .A(n1116), .Z(n18921) );
  BUF_X1 U1380 ( .A(n1114), .Z(n18924) );
  BUF_X1 U1381 ( .A(n1112), .Z(n18927) );
  BUF_X1 U1382 ( .A(n1110), .Z(n18930) );
  BUF_X1 U1383 ( .A(n1108), .Z(n18933) );
  BUF_X1 U1384 ( .A(n1106), .Z(n18936) );
  BUF_X1 U1385 ( .A(n1104), .Z(n18939) );
  BUF_X1 U1386 ( .A(n1102), .Z(n18942) );
  BUF_X1 U1387 ( .A(n1100), .Z(n18945) );
  BUF_X1 U1388 ( .A(n1098), .Z(n18948) );
  BUF_X1 U1389 ( .A(n1096), .Z(n18951) );
  BUF_X1 U1390 ( .A(n1094), .Z(n18954) );
  BUF_X1 U1391 ( .A(n1092), .Z(n18957) );
  BUF_X1 U1392 ( .A(n1090), .Z(n18960) );
  BUF_X1 U1393 ( .A(n1088), .Z(n18963) );
  BUF_X1 U1394 ( .A(n1086), .Z(n18966) );
  BUF_X1 U1395 ( .A(n1084), .Z(n18969) );
  BUF_X1 U1396 ( .A(n1082), .Z(n18972) );
  BUF_X1 U1397 ( .A(n1080), .Z(n18975) );
  BUF_X1 U1398 ( .A(n1078), .Z(n18978) );
  BUF_X1 U1399 ( .A(n1076), .Z(n18981) );
  BUF_X1 U1400 ( .A(n1073), .Z(n18993) );
  OAI22_X1 U1401 ( .A1(n18590), .A2(n18963), .B1(n18586), .B2(n17519), .ZN(
        n2944) );
  OAI22_X1 U1402 ( .A1(n18590), .A2(n18966), .B1(n18587), .B2(n17520), .ZN(
        n2945) );
  OAI22_X1 U1403 ( .A1(n18590), .A2(n18969), .B1(n18586), .B2(n17521), .ZN(
        n2946) );
  OAI22_X1 U1404 ( .A1(n18589), .A2(n18972), .B1(n18587), .B2(n17522), .ZN(
        n2947) );
  OAI22_X1 U1405 ( .A1(n18589), .A2(n18975), .B1(n18586), .B2(n17523), .ZN(
        n2948) );
  OAI22_X1 U1406 ( .A1(n18589), .A2(n18978), .B1(n18587), .B2(n17524), .ZN(
        n2949) );
  OAI22_X1 U1407 ( .A1(n18589), .A2(n18981), .B1(n18586), .B2(n17525), .ZN(
        n2950) );
  OAI22_X1 U1408 ( .A1(n18592), .A2(n18993), .B1(n18587), .B2(n17526), .ZN(
        n2951) );
  OAI22_X1 U1409 ( .A1(n18615), .A2(n18963), .B1(n2011), .B2(n17423), .ZN(
        n3008) );
  OAI22_X1 U1410 ( .A1(n18615), .A2(n18966), .B1(n18612), .B2(n17424), .ZN(
        n3009) );
  OAI22_X1 U1411 ( .A1(n18615), .A2(n18969), .B1(n18612), .B2(n17425), .ZN(
        n3010) );
  OAI22_X1 U1412 ( .A1(n18614), .A2(n18972), .B1(n18612), .B2(n17426), .ZN(
        n3011) );
  OAI22_X1 U1413 ( .A1(n18614), .A2(n18975), .B1(n18612), .B2(n17427), .ZN(
        n3012) );
  OAI22_X1 U1414 ( .A1(n18614), .A2(n18978), .B1(n18612), .B2(n17428), .ZN(
        n3013) );
  OAI22_X1 U1415 ( .A1(n18614), .A2(n18981), .B1(n18612), .B2(n17429), .ZN(
        n3014) );
  OAI22_X1 U1416 ( .A1(n18617), .A2(n18993), .B1(n2011), .B2(n17430), .ZN(
        n3015) );
  OAI22_X1 U1417 ( .A1(n18626), .A2(n18963), .B1(n1977), .B2(n17904), .ZN(
        n3040) );
  OAI22_X1 U1418 ( .A1(n18626), .A2(n18966), .B1(n18623), .B2(n17905), .ZN(
        n3041) );
  OAI22_X1 U1419 ( .A1(n18626), .A2(n18969), .B1(n18623), .B2(n17906), .ZN(
        n3042) );
  OAI22_X1 U1420 ( .A1(n18625), .A2(n18972), .B1(n18623), .B2(n17907), .ZN(
        n3043) );
  OAI22_X1 U1421 ( .A1(n18625), .A2(n18975), .B1(n18623), .B2(n17908), .ZN(
        n3044) );
  OAI22_X1 U1422 ( .A1(n18625), .A2(n18978), .B1(n18623), .B2(n17909), .ZN(
        n3045) );
  OAI22_X1 U1423 ( .A1(n18624), .A2(n18981), .B1(n18623), .B2(n17910), .ZN(
        n3046) );
  OAI22_X1 U1424 ( .A1(n18628), .A2(n18993), .B1(n1977), .B2(n17911), .ZN(
        n3047) );
  OAI22_X1 U1425 ( .A1(n18637), .A2(n18963), .B1(n1942), .B2(n17359), .ZN(
        n3072) );
  OAI22_X1 U1426 ( .A1(n18637), .A2(n18966), .B1(n18634), .B2(n17360), .ZN(
        n3073) );
  OAI22_X1 U1427 ( .A1(n18636), .A2(n18969), .B1(n18634), .B2(n17361), .ZN(
        n3074) );
  OAI22_X1 U1428 ( .A1(n18636), .A2(n18972), .B1(n18634), .B2(n17362), .ZN(
        n3075) );
  OAI22_X1 U1429 ( .A1(n18636), .A2(n18975), .B1(n18634), .B2(n17363), .ZN(
        n3076) );
  OAI22_X1 U1430 ( .A1(n18635), .A2(n18978), .B1(n18634), .B2(n17364), .ZN(
        n3077) );
  OAI22_X1 U1431 ( .A1(n18636), .A2(n18981), .B1(n18634), .B2(n17365), .ZN(
        n3078) );
  OAI22_X1 U1432 ( .A1(n18639), .A2(n18993), .B1(n1942), .B2(n17366), .ZN(
        n3079) );
  OAI22_X1 U1433 ( .A1(n18662), .A2(n18962), .B1(n1874), .B2(n17775), .ZN(
        n3136) );
  OAI22_X1 U1434 ( .A1(n18662), .A2(n18965), .B1(n18659), .B2(n17776), .ZN(
        n3137) );
  OAI22_X1 U1435 ( .A1(n18662), .A2(n18968), .B1(n18659), .B2(n17777), .ZN(
        n3138) );
  OAI22_X1 U1436 ( .A1(n18661), .A2(n18971), .B1(n18659), .B2(n17778), .ZN(
        n3139) );
  OAI22_X1 U1437 ( .A1(n18661), .A2(n18974), .B1(n18659), .B2(n17779), .ZN(
        n3140) );
  OAI22_X1 U1438 ( .A1(n18661), .A2(n18977), .B1(n18659), .B2(n17780), .ZN(
        n3141) );
  OAI22_X1 U1439 ( .A1(n18661), .A2(n18980), .B1(n18659), .B2(n17781), .ZN(
        n3142) );
  OAI22_X1 U1440 ( .A1(n18664), .A2(n18992), .B1(n1874), .B2(n17782), .ZN(
        n3143) );
  OAI22_X1 U1441 ( .A1(n18673), .A2(n18962), .B1(n1840), .B2(n17614), .ZN(
        n3168) );
  OAI22_X1 U1442 ( .A1(n18673), .A2(n18965), .B1(n18670), .B2(n17615), .ZN(
        n3169) );
  OAI22_X1 U1443 ( .A1(n18673), .A2(n18968), .B1(n18670), .B2(n17616), .ZN(
        n3170) );
  OAI22_X1 U1444 ( .A1(n18672), .A2(n18971), .B1(n18670), .B2(n17617), .ZN(
        n3171) );
  OAI22_X1 U1445 ( .A1(n18672), .A2(n18974), .B1(n18670), .B2(n17618), .ZN(
        n3172) );
  OAI22_X1 U1446 ( .A1(n18672), .A2(n18977), .B1(n18670), .B2(n17619), .ZN(
        n3173) );
  OAI22_X1 U1447 ( .A1(n18671), .A2(n18980), .B1(n18670), .B2(n17620), .ZN(
        n3174) );
  OAI22_X1 U1448 ( .A1(n18675), .A2(n18992), .B1(n1840), .B2(n17621), .ZN(
        n3175) );
  OAI22_X1 U1449 ( .A1(n18695), .A2(n18962), .B1(n1770), .B2(n18128), .ZN(
        n3232) );
  OAI22_X1 U1450 ( .A1(n18695), .A2(n18965), .B1(n18692), .B2(n18129), .ZN(
        n3233) );
  OAI22_X1 U1451 ( .A1(n18695), .A2(n18968), .B1(n18692), .B2(n18130), .ZN(
        n3234) );
  OAI22_X1 U1452 ( .A1(n18694), .A2(n18971), .B1(n18692), .B2(n18131), .ZN(
        n3235) );
  OAI22_X1 U1453 ( .A1(n18694), .A2(n18974), .B1(n18692), .B2(n18132), .ZN(
        n3236) );
  OAI22_X1 U1454 ( .A1(n18694), .A2(n18977), .B1(n18692), .B2(n18133), .ZN(
        n3237) );
  OAI22_X1 U1455 ( .A1(n18694), .A2(n18980), .B1(n18692), .B2(n18134), .ZN(
        n3238) );
  OAI22_X1 U1456 ( .A1(n18697), .A2(n18992), .B1(n1770), .B2(n18135), .ZN(
        n3239) );
  OAI22_X1 U1457 ( .A1(n18706), .A2(n18962), .B1(n1736), .B2(n17872), .ZN(
        n3264) );
  OAI22_X1 U1458 ( .A1(n18706), .A2(n18965), .B1(n18703), .B2(n17873), .ZN(
        n3265) );
  OAI22_X1 U1459 ( .A1(n18705), .A2(n18968), .B1(n18703), .B2(n17874), .ZN(
        n3266) );
  OAI22_X1 U1460 ( .A1(n18705), .A2(n18971), .B1(n18703), .B2(n17875), .ZN(
        n3267) );
  OAI22_X1 U1461 ( .A1(n18705), .A2(n18974), .B1(n18703), .B2(n17876), .ZN(
        n3268) );
  OAI22_X1 U1462 ( .A1(n18705), .A2(n18977), .B1(n18703), .B2(n17877), .ZN(
        n3269) );
  OAI22_X1 U1463 ( .A1(n18704), .A2(n18980), .B1(n18703), .B2(n17878), .ZN(
        n3270) );
  OAI22_X1 U1464 ( .A1(n18708), .A2(n18992), .B1(n1736), .B2(n17879), .ZN(
        n3271) );
  OAI22_X1 U1465 ( .A1(n18717), .A2(n18962), .B1(n1702), .B2(n17743), .ZN(
        n3296) );
  OAI22_X1 U1466 ( .A1(n18717), .A2(n18965), .B1(n18714), .B2(n17744), .ZN(
        n3297) );
  OAI22_X1 U1467 ( .A1(n18716), .A2(n18968), .B1(n18714), .B2(n17745), .ZN(
        n3298) );
  OAI22_X1 U1468 ( .A1(n18716), .A2(n18971), .B1(n18714), .B2(n17746), .ZN(
        n3299) );
  OAI22_X1 U1469 ( .A1(n18716), .A2(n18974), .B1(n18714), .B2(n17747), .ZN(
        n3300) );
  OAI22_X1 U1470 ( .A1(n18715), .A2(n18977), .B1(n18714), .B2(n17748), .ZN(
        n3301) );
  OAI22_X1 U1471 ( .A1(n18715), .A2(n18980), .B1(n18714), .B2(n17749), .ZN(
        n3302) );
  OAI22_X1 U1472 ( .A1(n18719), .A2(n18992), .B1(n1702), .B2(n17750), .ZN(
        n3303) );
  OAI22_X1 U1473 ( .A1(n18728), .A2(n18962), .B1(n1666), .B2(n18064), .ZN(
        n3328) );
  OAI22_X1 U1474 ( .A1(n18727), .A2(n18965), .B1(n18725), .B2(n18065), .ZN(
        n3329) );
  OAI22_X1 U1475 ( .A1(n18727), .A2(n18968), .B1(n18725), .B2(n18066), .ZN(
        n3330) );
  OAI22_X1 U1476 ( .A1(n18727), .A2(n18971), .B1(n18725), .B2(n18067), .ZN(
        n3331) );
  OAI22_X1 U1477 ( .A1(n18727), .A2(n18974), .B1(n18725), .B2(n18068), .ZN(
        n3332) );
  OAI22_X1 U1478 ( .A1(n18726), .A2(n18977), .B1(n18725), .B2(n18069), .ZN(
        n3333) );
  OAI22_X1 U1479 ( .A1(n18726), .A2(n18980), .B1(n18725), .B2(n18070), .ZN(
        n3334) );
  OAI22_X1 U1480 ( .A1(n18730), .A2(n18992), .B1(n1666), .B2(n18071), .ZN(
        n3335) );
  OAI22_X1 U1481 ( .A1(n18753), .A2(n18962), .B1(n18750), .B2(n17840), .ZN(
        n3392) );
  OAI22_X1 U1482 ( .A1(n18753), .A2(n18965), .B1(n18750), .B2(n17841), .ZN(
        n3393) );
  OAI22_X1 U1483 ( .A1(n18753), .A2(n18968), .B1(n18750), .B2(n17842), .ZN(
        n3394) );
  OAI22_X1 U1484 ( .A1(n18752), .A2(n18971), .B1(n1597), .B2(n17843), .ZN(
        n3395) );
  OAI22_X1 U1485 ( .A1(n18752), .A2(n18974), .B1(n18750), .B2(n17844), .ZN(
        n3396) );
  OAI22_X1 U1486 ( .A1(n18752), .A2(n18977), .B1(n1597), .B2(n17845), .ZN(
        n3397) );
  OAI22_X1 U1487 ( .A1(n18752), .A2(n18980), .B1(n18750), .B2(n17846), .ZN(
        n3398) );
  OAI22_X1 U1488 ( .A1(n18755), .A2(n18992), .B1(n1597), .B2(n17847), .ZN(
        n3399) );
  OAI22_X1 U1489 ( .A1(n18764), .A2(n18962), .B1(n18761), .B2(n18160), .ZN(
        n3424) );
  OAI22_X1 U1490 ( .A1(n18764), .A2(n18965), .B1(n18761), .B2(n18161), .ZN(
        n3425) );
  OAI22_X1 U1491 ( .A1(n18764), .A2(n18968), .B1(n18761), .B2(n18162), .ZN(
        n3426) );
  OAI22_X1 U1492 ( .A1(n18763), .A2(n18971), .B1(n1563), .B2(n18163), .ZN(
        n3427) );
  OAI22_X1 U1493 ( .A1(n18763), .A2(n18974), .B1(n18761), .B2(n18164), .ZN(
        n3428) );
  OAI22_X1 U1494 ( .A1(n18763), .A2(n18977), .B1(n1563), .B2(n18165), .ZN(
        n3429) );
  OAI22_X1 U1495 ( .A1(n18763), .A2(n18980), .B1(n18761), .B2(n18166), .ZN(
        n3430) );
  OAI22_X1 U1496 ( .A1(n18766), .A2(n18992), .B1(n1563), .B2(n18167), .ZN(
        n3431) );
  OAI22_X1 U1497 ( .A1(n18775), .A2(n18962), .B1(n18772), .B2(n18000), .ZN(
        n3456) );
  OAI22_X1 U1498 ( .A1(n18775), .A2(n18965), .B1(n18772), .B2(n18001), .ZN(
        n3457) );
  OAI22_X1 U1499 ( .A1(n18774), .A2(n18968), .B1(n18772), .B2(n18002), .ZN(
        n3458) );
  OAI22_X1 U1500 ( .A1(n18774), .A2(n18971), .B1(n1528), .B2(n18003), .ZN(
        n3459) );
  OAI22_X1 U1501 ( .A1(n18774), .A2(n18974), .B1(n18772), .B2(n18004), .ZN(
        n3460) );
  OAI22_X1 U1502 ( .A1(n18774), .A2(n18977), .B1(n1528), .B2(n18005), .ZN(
        n3461) );
  OAI22_X1 U1503 ( .A1(n18773), .A2(n18980), .B1(n18772), .B2(n18006), .ZN(
        n3462) );
  OAI22_X1 U1504 ( .A1(n18777), .A2(n18992), .B1(n1528), .B2(n18007), .ZN(
        n3463) );
  OAI22_X1 U1505 ( .A1(n18786), .A2(n18961), .B1(n18783), .B2(n18072), .ZN(
        n3488) );
  OAI22_X1 U1506 ( .A1(n18786), .A2(n18964), .B1(n18783), .B2(n18073), .ZN(
        n3489) );
  OAI22_X1 U1507 ( .A1(n18786), .A2(n18967), .B1(n18783), .B2(n18074), .ZN(
        n3490) );
  OAI22_X1 U1508 ( .A1(n18785), .A2(n18970), .B1(n1494), .B2(n18075), .ZN(
        n3491) );
  OAI22_X1 U1509 ( .A1(n18785), .A2(n18973), .B1(n18783), .B2(n18076), .ZN(
        n3492) );
  OAI22_X1 U1510 ( .A1(n18785), .A2(n18976), .B1(n1494), .B2(n18077), .ZN(
        n3493) );
  OAI22_X1 U1511 ( .A1(n18785), .A2(n18979), .B1(n18783), .B2(n18078), .ZN(
        n3494) );
  OAI22_X1 U1512 ( .A1(n18788), .A2(n18991), .B1(n1494), .B2(n18079), .ZN(
        n3495) );
  OAI22_X1 U1513 ( .A1(n18797), .A2(n18961), .B1(n18794), .B2(n17527), .ZN(
        n3520) );
  OAI22_X1 U1514 ( .A1(n18797), .A2(n18964), .B1(n18794), .B2(n17528), .ZN(
        n3521) );
  OAI22_X1 U1515 ( .A1(n18796), .A2(n18967), .B1(n18794), .B2(n17529), .ZN(
        n3522) );
  OAI22_X1 U1516 ( .A1(n18796), .A2(n18970), .B1(n1460), .B2(n17530), .ZN(
        n3523) );
  OAI22_X1 U1517 ( .A1(n18796), .A2(n18973), .B1(n18794), .B2(n17531), .ZN(
        n3524) );
  OAI22_X1 U1518 ( .A1(n18796), .A2(n18976), .B1(n1460), .B2(n17532), .ZN(
        n3525) );
  OAI22_X1 U1519 ( .A1(n18795), .A2(n18979), .B1(n18794), .B2(n17533), .ZN(
        n3526) );
  OAI22_X1 U1520 ( .A1(n18799), .A2(n18991), .B1(n1460), .B2(n17534), .ZN(
        n3527) );
  OAI22_X1 U1521 ( .A1(n18808), .A2(n18961), .B1(n18805), .B2(n17391), .ZN(
        n3552) );
  OAI22_X1 U1522 ( .A1(n18808), .A2(n18964), .B1(n18805), .B2(n17392), .ZN(
        n3553) );
  OAI22_X1 U1523 ( .A1(n18807), .A2(n18967), .B1(n18805), .B2(n17393), .ZN(
        n3554) );
  OAI22_X1 U1524 ( .A1(n18807), .A2(n18970), .B1(n1426), .B2(n17394), .ZN(
        n3555) );
  OAI22_X1 U1525 ( .A1(n18807), .A2(n18973), .B1(n18805), .B2(n17395), .ZN(
        n3556) );
  OAI22_X1 U1526 ( .A1(n18807), .A2(n18976), .B1(n1426), .B2(n17396), .ZN(
        n3557) );
  OAI22_X1 U1527 ( .A1(n18806), .A2(n18979), .B1(n18805), .B2(n17397), .ZN(
        n3558) );
  OAI22_X1 U1528 ( .A1(n18810), .A2(n18991), .B1(n1426), .B2(n17398), .ZN(
        n3559) );
  OAI22_X1 U1529 ( .A1(n18819), .A2(n18961), .B1(n18816), .B2(n17679), .ZN(
        n3584) );
  OAI22_X1 U1530 ( .A1(n18818), .A2(n18964), .B1(n18816), .B2(n17680), .ZN(
        n3585) );
  OAI22_X1 U1531 ( .A1(n18818), .A2(n18967), .B1(n18816), .B2(n17681), .ZN(
        n3586) );
  OAI22_X1 U1532 ( .A1(n18818), .A2(n18970), .B1(n1390), .B2(n17682), .ZN(
        n3587) );
  OAI22_X1 U1533 ( .A1(n18818), .A2(n18973), .B1(n18816), .B2(n17683), .ZN(
        n3588) );
  OAI22_X1 U1534 ( .A1(n18817), .A2(n18976), .B1(n1390), .B2(n17684), .ZN(
        n3589) );
  OAI22_X1 U1535 ( .A1(n18817), .A2(n18979), .B1(n18816), .B2(n17685), .ZN(
        n3590) );
  OAI22_X1 U1536 ( .A1(n18821), .A2(n18991), .B1(n1390), .B2(n17686), .ZN(
        n3591) );
  OAI22_X1 U1537 ( .A1(n18834), .A2(n18961), .B1(n18827), .B2(n17807), .ZN(
        n3616) );
  OAI22_X1 U1538 ( .A1(n18834), .A2(n18964), .B1(n18827), .B2(n17808), .ZN(
        n3617) );
  OAI22_X1 U1539 ( .A1(n18834), .A2(n18967), .B1(n18827), .B2(n17809), .ZN(
        n3618) );
  OAI22_X1 U1540 ( .A1(n18834), .A2(n18970), .B1(n1356), .B2(n17810), .ZN(
        n3619) );
  OAI22_X1 U1541 ( .A1(n18835), .A2(n18973), .B1(n18827), .B2(n17811), .ZN(
        n3620) );
  OAI22_X1 U1542 ( .A1(n18835), .A2(n18976), .B1(n1356), .B2(n17812), .ZN(
        n3621) );
  OAI22_X1 U1543 ( .A1(n18835), .A2(n18979), .B1(n18827), .B2(n17813), .ZN(
        n3622) );
  OAI22_X1 U1544 ( .A1(n18835), .A2(n18991), .B1(n1356), .B2(n17814), .ZN(
        n3623) );
  OAI22_X1 U1545 ( .A1(n18841), .A2(n18961), .B1(n18838), .B2(n17327), .ZN(
        n3648) );
  OAI22_X1 U1546 ( .A1(n18841), .A2(n18964), .B1(n18838), .B2(n17328), .ZN(
        n3649) );
  OAI22_X1 U1547 ( .A1(n18840), .A2(n18967), .B1(n18838), .B2(n17329), .ZN(
        n3650) );
  OAI22_X1 U1548 ( .A1(n18840), .A2(n18970), .B1(n1322), .B2(n17330), .ZN(
        n3651) );
  OAI22_X1 U1549 ( .A1(n18840), .A2(n18973), .B1(n18838), .B2(n17331), .ZN(
        n3652) );
  OAI22_X1 U1550 ( .A1(n18840), .A2(n18976), .B1(n1322), .B2(n17332), .ZN(
        n3653) );
  OAI22_X1 U1551 ( .A1(n18839), .A2(n18979), .B1(n18838), .B2(n17333), .ZN(
        n3654) );
  OAI22_X1 U1552 ( .A1(n18843), .A2(n18991), .B1(n1322), .B2(n17334), .ZN(
        n3655) );
  OAI22_X1 U1553 ( .A1(n18852), .A2(n18961), .B1(n18849), .B2(n18008), .ZN(
        n3680) );
  OAI22_X1 U1554 ( .A1(n18852), .A2(n18964), .B1(n18849), .B2(n18009), .ZN(
        n3681) );
  OAI22_X1 U1555 ( .A1(n18851), .A2(n18967), .B1(n18849), .B2(n18010), .ZN(
        n3682) );
  OAI22_X1 U1556 ( .A1(n18851), .A2(n18970), .B1(n1288), .B2(n18011), .ZN(
        n3683) );
  OAI22_X1 U1557 ( .A1(n18851), .A2(n18973), .B1(n18849), .B2(n18012), .ZN(
        n3684) );
  OAI22_X1 U1558 ( .A1(n18851), .A2(n18976), .B1(n1288), .B2(n18013), .ZN(
        n3685) );
  OAI22_X1 U1559 ( .A1(n18850), .A2(n18979), .B1(n18849), .B2(n18014), .ZN(
        n3686) );
  OAI22_X1 U1560 ( .A1(n18854), .A2(n18991), .B1(n1288), .B2(n18015), .ZN(
        n3687) );
  OAI22_X1 U1561 ( .A1(n18863), .A2(n18961), .B1(n18860), .B2(n18254), .ZN(
        n3712) );
  OAI22_X1 U1562 ( .A1(n18862), .A2(n18964), .B1(n18860), .B2(n18255), .ZN(
        n3713) );
  OAI22_X1 U1563 ( .A1(n18862), .A2(n18967), .B1(n18860), .B2(n18256), .ZN(
        n3714) );
  OAI22_X1 U1564 ( .A1(n18862), .A2(n18970), .B1(n1252), .B2(n18257), .ZN(
        n3715) );
  OAI22_X1 U1565 ( .A1(n18862), .A2(n18973), .B1(n18860), .B2(n18258), .ZN(
        n3716) );
  OAI22_X1 U1566 ( .A1(n18861), .A2(n18976), .B1(n1252), .B2(n18259), .ZN(
        n3717) );
  OAI22_X1 U1567 ( .A1(n18861), .A2(n18979), .B1(n18860), .B2(n18260), .ZN(
        n3718) );
  OAI22_X1 U1568 ( .A1(n18865), .A2(n18991), .B1(n1252), .B2(n18261), .ZN(
        n3719) );
  OAI22_X1 U1569 ( .A1(n18878), .A2(n18961), .B1(n18871), .B2(n17968), .ZN(
        n3744) );
  OAI22_X1 U1570 ( .A1(n18878), .A2(n18964), .B1(n1214), .B2(n17969), .ZN(
        n3745) );
  OAI22_X1 U1571 ( .A1(n18878), .A2(n18967), .B1(n18871), .B2(n17970), .ZN(
        n3746) );
  OAI22_X1 U1572 ( .A1(n18878), .A2(n18970), .B1(n1214), .B2(n17971), .ZN(
        n3747) );
  OAI22_X1 U1573 ( .A1(n18879), .A2(n18973), .B1(n18871), .B2(n17972), .ZN(
        n3748) );
  OAI22_X1 U1574 ( .A1(n18879), .A2(n18976), .B1(n1214), .B2(n17973), .ZN(
        n3749) );
  OAI22_X1 U1575 ( .A1(n18879), .A2(n18979), .B1(n18871), .B2(n17974), .ZN(
        n3750) );
  OAI22_X1 U1576 ( .A1(n18879), .A2(n18991), .B1(n1214), .B2(n17975), .ZN(
        n3751) );
  OAI22_X1 U1577 ( .A1(n18885), .A2(n18961), .B1(n18882), .B2(n17455), .ZN(
        n3776) );
  OAI22_X1 U1578 ( .A1(n18884), .A2(n18964), .B1(n1178), .B2(n17456), .ZN(
        n3777) );
  OAI22_X1 U1579 ( .A1(n18884), .A2(n18967), .B1(n18882), .B2(n17457), .ZN(
        n3778) );
  OAI22_X1 U1580 ( .A1(n18884), .A2(n18970), .B1(n1178), .B2(n17458), .ZN(
        n3779) );
  OAI22_X1 U1581 ( .A1(n18884), .A2(n18973), .B1(n18882), .B2(n17459), .ZN(
        n3780) );
  OAI22_X1 U1582 ( .A1(n18883), .A2(n18976), .B1(n1178), .B2(n17460), .ZN(
        n3781) );
  OAI22_X1 U1583 ( .A1(n18883), .A2(n18979), .B1(n18882), .B2(n17461), .ZN(
        n3782) );
  OAI22_X1 U1584 ( .A1(n18887), .A2(n18991), .B1(n1178), .B2(n17462), .ZN(
        n3783) );
  OAI22_X1 U1585 ( .A1(n18900), .A2(n18961), .B1(n18893), .B2(n17719), .ZN(
        n3808) );
  OAI22_X1 U1586 ( .A1(n18900), .A2(n18964), .B1(n1142), .B2(n17720), .ZN(
        n3809) );
  OAI22_X1 U1587 ( .A1(n18900), .A2(n18967), .B1(n18893), .B2(n17721), .ZN(
        n3810) );
  OAI22_X1 U1588 ( .A1(n18900), .A2(n18970), .B1(n1142), .B2(n17722), .ZN(
        n3811) );
  OAI22_X1 U1589 ( .A1(n18901), .A2(n18973), .B1(n18893), .B2(n17723), .ZN(
        n3812) );
  OAI22_X1 U1590 ( .A1(n18901), .A2(n18976), .B1(n1142), .B2(n17724), .ZN(
        n3813) );
  OAI22_X1 U1591 ( .A1(n18901), .A2(n18979), .B1(n18893), .B2(n17725), .ZN(
        n3814) );
  OAI22_X1 U1592 ( .A1(n18901), .A2(n18991), .B1(n1142), .B2(n17726), .ZN(
        n3815) );
  OAI22_X1 U1593 ( .A1(n18987), .A2(n18961), .B1(n1074), .B2(n17936), .ZN(
        n3840) );
  OAI22_X1 U1594 ( .A1(n18988), .A2(n18964), .B1(n1074), .B2(n17937), .ZN(
        n3841) );
  OAI22_X1 U1595 ( .A1(n18988), .A2(n18967), .B1(n1074), .B2(n17938), .ZN(
        n3842) );
  OAI22_X1 U1596 ( .A1(n18988), .A2(n18970), .B1(n1074), .B2(n17939), .ZN(
        n3843) );
  OAI22_X1 U1597 ( .A1(n18988), .A2(n18973), .B1(n1074), .B2(n17940), .ZN(
        n3844) );
  OAI22_X1 U1598 ( .A1(n18988), .A2(n18976), .B1(n18982), .B2(n17941), .ZN(
        n3845) );
  OAI22_X1 U1599 ( .A1(n18989), .A2(n18979), .B1(n18982), .B2(n17942), .ZN(
        n3846) );
  OAI22_X1 U1600 ( .A1(n18989), .A2(n18991), .B1(n1074), .B2(n17943), .ZN(
        n3847) );
  OAI22_X1 U1601 ( .A1(n18588), .A2(n1136), .B1(n18586), .B2(n17535), .ZN(
        n2920) );
  OAI22_X1 U1602 ( .A1(n18595), .A2(n1134), .B1(n18586), .B2(n17536), .ZN(
        n2921) );
  OAI22_X1 U1603 ( .A1(n18613), .A2(n1136), .B1(n18612), .B2(n17431), .ZN(
        n2984) );
  OAI22_X1 U1604 ( .A1(n18620), .A2(n1132), .B1(n18612), .B2(n17432), .ZN(
        n2986) );
  OAI22_X1 U1605 ( .A1(n18625), .A2(n1134), .B1(n18623), .B2(n17912), .ZN(
        n3017) );
  OAI22_X1 U1606 ( .A1(n18631), .A2(n1132), .B1(n18623), .B2(n17913), .ZN(
        n3018) );
  OAI22_X1 U1607 ( .A1(n18635), .A2(n1136), .B1(n18634), .B2(n17383), .ZN(
        n3048) );
  OAI22_X1 U1608 ( .A1(n18642), .A2(n1134), .B1(n18634), .B2(n17384), .ZN(
        n3049) );
  OAI22_X1 U1609 ( .A1(n18642), .A2(n1132), .B1(n18634), .B2(n17385), .ZN(
        n3050) );
  OAI22_X1 U1610 ( .A1(n18660), .A2(n1136), .B1(n18659), .B2(n17783), .ZN(
        n3112) );
  OAI22_X1 U1611 ( .A1(n18667), .A2(n1130), .B1(n18659), .B2(n17784), .ZN(
        n3115) );
  OAI22_X1 U1612 ( .A1(n18672), .A2(n1134), .B1(n18670), .B2(n17670), .ZN(
        n3145) );
  OAI22_X1 U1613 ( .A1(n18678), .A2(n1130), .B1(n18670), .B2(n17672), .ZN(
        n3147) );
  OAI22_X1 U1614 ( .A1(n18693), .A2(n1132), .B1(n18692), .B2(n18136), .ZN(
        n3210) );
  OAI22_X1 U1615 ( .A1(n18700), .A2(n1130), .B1(n18692), .B2(n18137), .ZN(
        n3211) );
  OAI22_X1 U1616 ( .A1(n18704), .A2(n1136), .B1(n18703), .B2(n17880), .ZN(
        n3240) );
  OAI22_X1 U1617 ( .A1(n18711), .A2(n1132), .B1(n18703), .B2(n17881), .ZN(
        n3242) );
  OAI22_X1 U1618 ( .A1(n18711), .A2(n1130), .B1(n18703), .B2(n17882), .ZN(
        n3243) );
  OAI22_X1 U1619 ( .A1(n18716), .A2(n1134), .B1(n18714), .B2(n17751), .ZN(
        n3273) );
  OAI22_X1 U1620 ( .A1(n18722), .A2(n1132), .B1(n18714), .B2(n17752), .ZN(
        n3274) );
  OAI22_X1 U1621 ( .A1(n18722), .A2(n1130), .B1(n18714), .B2(n17753), .ZN(
        n3275) );
  OAI22_X1 U1622 ( .A1(n18726), .A2(n1136), .B1(n18725), .B2(n18080), .ZN(
        n3304) );
  OAI22_X1 U1623 ( .A1(n18733), .A2(n1134), .B1(n18725), .B2(n18081), .ZN(
        n3305) );
  OAI22_X1 U1624 ( .A1(n18733), .A2(n1132), .B1(n18725), .B2(n18082), .ZN(
        n3306) );
  OAI22_X1 U1625 ( .A1(n18733), .A2(n1130), .B1(n18725), .B2(n18083), .ZN(
        n3307) );
  OAI22_X1 U1626 ( .A1(n18751), .A2(n1136), .B1(n18750), .B2(n17848), .ZN(
        n3368) );
  OAI22_X1 U1627 ( .A1(n18758), .A2(n1128), .B1(n18750), .B2(n17852), .ZN(
        n3372) );
  OAI22_X1 U1628 ( .A1(n18762), .A2(n1134), .B1(n18761), .B2(n18168), .ZN(
        n3401) );
  OAI22_X1 U1629 ( .A1(n18769), .A2(n1128), .B1(n18761), .B2(n18169), .ZN(
        n3404) );
  OAI22_X1 U1630 ( .A1(n18773), .A2(n1136), .B1(n18772), .B2(n18016), .ZN(
        n3432) );
  OAI22_X1 U1631 ( .A1(n18780), .A2(n1134), .B1(n18772), .B2(n18017), .ZN(
        n3433) );
  OAI22_X1 U1632 ( .A1(n18780), .A2(n1128), .B1(n18772), .B2(n18018), .ZN(
        n3436) );
  OAI22_X1 U1633 ( .A1(n18784), .A2(n1132), .B1(n18783), .B2(n18084), .ZN(
        n3466) );
  OAI22_X1 U1634 ( .A1(n18791), .A2(n1128), .B1(n18783), .B2(n18085), .ZN(
        n3468) );
  OAI22_X1 U1635 ( .A1(n18795), .A2(n1136), .B1(n18794), .B2(n17537), .ZN(
        n3496) );
  OAI22_X1 U1636 ( .A1(n18802), .A2(n1132), .B1(n18794), .B2(n17538), .ZN(
        n3498) );
  OAI22_X1 U1637 ( .A1(n18802), .A2(n1128), .B1(n18794), .B2(n17539), .ZN(
        n3500) );
  OAI22_X1 U1638 ( .A1(n18806), .A2(n1134), .B1(n18805), .B2(n17399), .ZN(
        n3529) );
  OAI22_X1 U1639 ( .A1(n18813), .A2(n1132), .B1(n18805), .B2(n17400), .ZN(
        n3530) );
  OAI22_X1 U1640 ( .A1(n18813), .A2(n1128), .B1(n18805), .B2(n17401), .ZN(
        n3532) );
  OAI22_X1 U1641 ( .A1(n18817), .A2(n1136), .B1(n18816), .B2(n17687), .ZN(
        n3560) );
  OAI22_X1 U1642 ( .A1(n18824), .A2(n1134), .B1(n18816), .B2(n17688), .ZN(
        n3561) );
  OAI22_X1 U1643 ( .A1(n18824), .A2(n1132), .B1(n18816), .B2(n17689), .ZN(
        n3562) );
  OAI22_X1 U1644 ( .A1(n18824), .A2(n1128), .B1(n18816), .B2(n17690), .ZN(
        n3564) );
  OAI22_X1 U1645 ( .A1(n18828), .A2(n1130), .B1(n18827), .B2(n17815), .ZN(
        n3595) );
  OAI22_X1 U1646 ( .A1(n18829), .A2(n1128), .B1(n18827), .B2(n17816), .ZN(
        n3596) );
  OAI22_X1 U1647 ( .A1(n18839), .A2(n1136), .B1(n18838), .B2(n17335), .ZN(
        n3624) );
  OAI22_X1 U1648 ( .A1(n18846), .A2(n1130), .B1(n18838), .B2(n17336), .ZN(
        n3627) );
  OAI22_X1 U1649 ( .A1(n18846), .A2(n1128), .B1(n18838), .B2(n17337), .ZN(
        n3628) );
  OAI22_X1 U1650 ( .A1(n18850), .A2(n1134), .B1(n18849), .B2(n18019), .ZN(
        n3657) );
  OAI22_X1 U1651 ( .A1(n18857), .A2(n1130), .B1(n18849), .B2(n18020), .ZN(
        n3659) );
  OAI22_X1 U1652 ( .A1(n18857), .A2(n1128), .B1(n18849), .B2(n18021), .ZN(
        n3660) );
  OAI22_X1 U1653 ( .A1(n18861), .A2(n1136), .B1(n18860), .B2(n18262), .ZN(
        n3688) );
  OAI22_X1 U1654 ( .A1(n18868), .A2(n1134), .B1(n18860), .B2(n18263), .ZN(
        n3689) );
  OAI22_X1 U1655 ( .A1(n18868), .A2(n1130), .B1(n18860), .B2(n18264), .ZN(
        n3691) );
  OAI22_X1 U1656 ( .A1(n18868), .A2(n1128), .B1(n18860), .B2(n18265), .ZN(
        n3692) );
  OAI22_X1 U1657 ( .A1(n18872), .A2(n1132), .B1(n18871), .B2(n17976), .ZN(
        n3722) );
  OAI22_X1 U1658 ( .A1(n18872), .A2(n1130), .B1(n18871), .B2(n17977), .ZN(
        n3723) );
  OAI22_X1 U1659 ( .A1(n18873), .A2(n1128), .B1(n18871), .B2(n17978), .ZN(
        n3724) );
  OAI22_X1 U1660 ( .A1(n18883), .A2(n1136), .B1(n18882), .B2(n17463), .ZN(
        n3752) );
  OAI22_X1 U1661 ( .A1(n18890), .A2(n1132), .B1(n18882), .B2(n17464), .ZN(
        n3754) );
  OAI22_X1 U1662 ( .A1(n18890), .A2(n1130), .B1(n18882), .B2(n17465), .ZN(
        n3755) );
  OAI22_X1 U1663 ( .A1(n18890), .A2(n1128), .B1(n18882), .B2(n17466), .ZN(
        n3756) );
  OAI22_X1 U1664 ( .A1(n18894), .A2(n1134), .B1(n18893), .B2(n17711), .ZN(
        n3785) );
  OAI22_X1 U1665 ( .A1(n18894), .A2(n1132), .B1(n18893), .B2(n17712), .ZN(
        n3786) );
  OAI22_X1 U1666 ( .A1(n18894), .A2(n1130), .B1(n18893), .B2(n17713), .ZN(
        n3787) );
  OAI22_X1 U1667 ( .A1(n18895), .A2(n1128), .B1(n18893), .B2(n17714), .ZN(
        n3788) );
  OAI22_X1 U1668 ( .A1(n18983), .A2(n1136), .B1(n18982), .B2(n17944), .ZN(
        n3816) );
  OAI22_X1 U1669 ( .A1(n18983), .A2(n1134), .B1(n18982), .B2(n17945), .ZN(
        n3817) );
  OAI22_X1 U1670 ( .A1(n18983), .A2(n1132), .B1(n18982), .B2(n17946), .ZN(
        n3818) );
  OAI22_X1 U1671 ( .A1(n18983), .A2(n1130), .B1(n18982), .B2(n17947), .ZN(
        n3819) );
  OAI22_X1 U1672 ( .A1(n18983), .A2(n1128), .B1(n18982), .B2(n17948), .ZN(
        n3820) );
  OAI22_X1 U1673 ( .A1(n18984), .A2(n18904), .B1(n18982), .B2(n17949), .ZN(
        n3821) );
  OAI22_X1 U1674 ( .A1(n18984), .A2(n18907), .B1(n18982), .B2(n17950), .ZN(
        n3822) );
  OAI22_X1 U1675 ( .A1(n18984), .A2(n18910), .B1(n18982), .B2(n17951), .ZN(
        n3823) );
  OAI22_X1 U1676 ( .A1(n18984), .A2(n18913), .B1(n18982), .B2(n17952), .ZN(
        n3824) );
  OAI22_X1 U1677 ( .A1(n18984), .A2(n18916), .B1(n18982), .B2(n17953), .ZN(
        n3825) );
  OAI22_X1 U1678 ( .A1(n18985), .A2(n18919), .B1(n18982), .B2(n17954), .ZN(
        n3826) );
  OAI22_X1 U1679 ( .A1(n18985), .A2(n18922), .B1(n18982), .B2(n17955), .ZN(
        n3827) );
  OAI22_X1 U1680 ( .A1(n18985), .A2(n18925), .B1(n18982), .B2(n17956), .ZN(
        n3828) );
  OAI22_X1 U1681 ( .A1(n18985), .A2(n18928), .B1(n18982), .B2(n17957), .ZN(
        n3829) );
  OAI22_X1 U1682 ( .A1(n18985), .A2(n18931), .B1(n18982), .B2(n17958), .ZN(
        n3830) );
  OAI22_X1 U1683 ( .A1(n18986), .A2(n18934), .B1(n1074), .B2(n17959), .ZN(
        n3831) );
  OAI22_X1 U1684 ( .A1(n18986), .A2(n18937), .B1(n1074), .B2(n17960), .ZN(
        n3832) );
  OAI22_X1 U1685 ( .A1(n18986), .A2(n18940), .B1(n1074), .B2(n17961), .ZN(
        n3833) );
  OAI22_X1 U1686 ( .A1(n18986), .A2(n18943), .B1(n1074), .B2(n17962), .ZN(
        n3834) );
  OAI22_X1 U1687 ( .A1(n18986), .A2(n18946), .B1(n1074), .B2(n17963), .ZN(
        n3835) );
  OAI22_X1 U1688 ( .A1(n18987), .A2(n18949), .B1(n18982), .B2(n17964), .ZN(
        n3836) );
  OAI22_X1 U1689 ( .A1(n18987), .A2(n18952), .B1(n18982), .B2(n17965), .ZN(
        n3837) );
  OAI22_X1 U1690 ( .A1(n18987), .A2(n18955), .B1(n18982), .B2(n17966), .ZN(
        n3838) );
  OAI22_X1 U1691 ( .A1(n18987), .A2(n18958), .B1(n18982), .B2(n17967), .ZN(
        n3839) );
  OAI22_X1 U1692 ( .A1(n1282), .A2(n18588), .B1(n18586), .B2(n17540), .ZN(
        n2922) );
  OAI22_X1 U1693 ( .A1(n1419), .A2(n18588), .B1(n18586), .B2(n17541), .ZN(
        n2923) );
  OAI22_X1 U1694 ( .A1(n1694), .A2(n18588), .B1(n18586), .B2(n17542), .ZN(
        n2924) );
  OAI22_X1 U1695 ( .A1(n18595), .A2(n18906), .B1(n18586), .B2(n17543), .ZN(
        n2925) );
  OAI22_X1 U1696 ( .A1(n18595), .A2(n18909), .B1(n18586), .B2(n17544), .ZN(
        n2926) );
  OAI22_X1 U1697 ( .A1(n18595), .A2(n18912), .B1(n18586), .B2(n17545), .ZN(
        n2927) );
  OAI22_X1 U1698 ( .A1(n18594), .A2(n18915), .B1(n18586), .B2(n17546), .ZN(
        n2928) );
  OAI22_X1 U1699 ( .A1(n18594), .A2(n18918), .B1(n18586), .B2(n17547), .ZN(
        n2929) );
  OAI22_X1 U1700 ( .A1(n18594), .A2(n18921), .B1(n18586), .B2(n17548), .ZN(
        n2930) );
  OAI22_X1 U1701 ( .A1(n18594), .A2(n18924), .B1(n18586), .B2(n17549), .ZN(
        n2931) );
  OAI22_X1 U1702 ( .A1(n18593), .A2(n18927), .B1(n18587), .B2(n17550), .ZN(
        n2932) );
  OAI22_X1 U1703 ( .A1(n18593), .A2(n18930), .B1(n18587), .B2(n17551), .ZN(
        n2933) );
  OAI22_X1 U1704 ( .A1(n18593), .A2(n18933), .B1(n18587), .B2(n17552), .ZN(
        n2934) );
  OAI22_X1 U1705 ( .A1(n18593), .A2(n18936), .B1(n18587), .B2(n17553), .ZN(
        n2935) );
  OAI22_X1 U1706 ( .A1(n18592), .A2(n18939), .B1(n18587), .B2(n17554), .ZN(
        n2936) );
  OAI22_X1 U1707 ( .A1(n18592), .A2(n18942), .B1(n18587), .B2(n17555), .ZN(
        n2937) );
  OAI22_X1 U1708 ( .A1(n18592), .A2(n18945), .B1(n18587), .B2(n17556), .ZN(
        n2938) );
  OAI22_X1 U1709 ( .A1(n18591), .A2(n18948), .B1(n18587), .B2(n17557), .ZN(
        n2939) );
  OAI22_X1 U1710 ( .A1(n18591), .A2(n18951), .B1(n18587), .B2(n17558), .ZN(
        n2940) );
  OAI22_X1 U1711 ( .A1(n18591), .A2(n18954), .B1(n18587), .B2(n17559), .ZN(
        n2941) );
  OAI22_X1 U1712 ( .A1(n18591), .A2(n18957), .B1(n18587), .B2(n17560), .ZN(
        n2942) );
  OAI22_X1 U1713 ( .A1(n18590), .A2(n18960), .B1(n18587), .B2(n17561), .ZN(
        n2943) );
  OAI22_X1 U1714 ( .A1(n1209), .A2(n18613), .B1(n18612), .B2(n17433), .ZN(
        n2985) );
  OAI22_X1 U1715 ( .A1(n1419), .A2(n18613), .B1(n18612), .B2(n17434), .ZN(
        n2987) );
  OAI22_X1 U1716 ( .A1(n1694), .A2(n18613), .B1(n18612), .B2(n17435), .ZN(
        n2988) );
  OAI22_X1 U1717 ( .A1(n18620), .A2(n18906), .B1(n18612), .B2(n17436), .ZN(
        n2989) );
  OAI22_X1 U1718 ( .A1(n18620), .A2(n18909), .B1(n18612), .B2(n17437), .ZN(
        n2990) );
  OAI22_X1 U1719 ( .A1(n18620), .A2(n18912), .B1(n18612), .B2(n17438), .ZN(
        n2991) );
  OAI22_X1 U1720 ( .A1(n18619), .A2(n18915), .B1(n18612), .B2(n17439), .ZN(
        n2992) );
  OAI22_X1 U1721 ( .A1(n18619), .A2(n18918), .B1(n18612), .B2(n17440), .ZN(
        n2993) );
  OAI22_X1 U1722 ( .A1(n18619), .A2(n18921), .B1(n18612), .B2(n17441), .ZN(
        n2994) );
  OAI22_X1 U1723 ( .A1(n18619), .A2(n18924), .B1(n18612), .B2(n17442), .ZN(
        n2995) );
  OAI22_X1 U1724 ( .A1(n18618), .A2(n18927), .B1(n2011), .B2(n17443), .ZN(
        n2996) );
  OAI22_X1 U1725 ( .A1(n18618), .A2(n18930), .B1(n2011), .B2(n17444), .ZN(
        n2997) );
  OAI22_X1 U1726 ( .A1(n18618), .A2(n18933), .B1(n2011), .B2(n17445), .ZN(
        n2998) );
  OAI22_X1 U1727 ( .A1(n18618), .A2(n18936), .B1(n2011), .B2(n17446), .ZN(
        n2999) );
  OAI22_X1 U1728 ( .A1(n18617), .A2(n18939), .B1(n2011), .B2(n17447), .ZN(
        n3000) );
  OAI22_X1 U1729 ( .A1(n18617), .A2(n18942), .B1(n2011), .B2(n17448), .ZN(
        n3001) );
  OAI22_X1 U1730 ( .A1(n18617), .A2(n18945), .B1(n2011), .B2(n17449), .ZN(
        n3002) );
  OAI22_X1 U1731 ( .A1(n18616), .A2(n18948), .B1(n2011), .B2(n17450), .ZN(
        n3003) );
  OAI22_X1 U1732 ( .A1(n18616), .A2(n18951), .B1(n2011), .B2(n17451), .ZN(
        n3004) );
  OAI22_X1 U1733 ( .A1(n18616), .A2(n18954), .B1(n18612), .B2(n17452), .ZN(
        n3005) );
  OAI22_X1 U1734 ( .A1(n18616), .A2(n18957), .B1(n18612), .B2(n17453), .ZN(
        n3006) );
  OAI22_X1 U1735 ( .A1(n18615), .A2(n18960), .B1(n18612), .B2(n17454), .ZN(
        n3007) );
  OAI22_X1 U1736 ( .A1(n1174), .A2(n18624), .B1(n18623), .B2(n17914), .ZN(
        n3016) );
  OAI22_X1 U1737 ( .A1(n1419), .A2(n18624), .B1(n18623), .B2(n17915), .ZN(
        n3019) );
  OAI22_X1 U1738 ( .A1(n1694), .A2(n18624), .B1(n18623), .B2(n17916), .ZN(
        n3020) );
  OAI22_X1 U1739 ( .A1(n18631), .A2(n18906), .B1(n18623), .B2(n17917), .ZN(
        n3021) );
  OAI22_X1 U1740 ( .A1(n18631), .A2(n18909), .B1(n18623), .B2(n17918), .ZN(
        n3022) );
  OAI22_X1 U1741 ( .A1(n18631), .A2(n18912), .B1(n18623), .B2(n17919), .ZN(
        n3023) );
  OAI22_X1 U1742 ( .A1(n18630), .A2(n18915), .B1(n18623), .B2(n17920), .ZN(
        n3024) );
  OAI22_X1 U1743 ( .A1(n18630), .A2(n18918), .B1(n18623), .B2(n17921), .ZN(
        n3025) );
  OAI22_X1 U1744 ( .A1(n18630), .A2(n18921), .B1(n18623), .B2(n17922), .ZN(
        n3026) );
  OAI22_X1 U1745 ( .A1(n18630), .A2(n18924), .B1(n18623), .B2(n17923), .ZN(
        n3027) );
  OAI22_X1 U1746 ( .A1(n18629), .A2(n18927), .B1(n1977), .B2(n17924), .ZN(
        n3028) );
  OAI22_X1 U1747 ( .A1(n18629), .A2(n18930), .B1(n1977), .B2(n17925), .ZN(
        n3029) );
  OAI22_X1 U1748 ( .A1(n18629), .A2(n18933), .B1(n1977), .B2(n17926), .ZN(
        n3030) );
  OAI22_X1 U1749 ( .A1(n18629), .A2(n18936), .B1(n1977), .B2(n17927), .ZN(
        n3031) );
  OAI22_X1 U1750 ( .A1(n18628), .A2(n18939), .B1(n1977), .B2(n17928), .ZN(
        n3032) );
  OAI22_X1 U1751 ( .A1(n18628), .A2(n18942), .B1(n1977), .B2(n17929), .ZN(
        n3033) );
  OAI22_X1 U1752 ( .A1(n18628), .A2(n18945), .B1(n1977), .B2(n17930), .ZN(
        n3034) );
  OAI22_X1 U1753 ( .A1(n18627), .A2(n18948), .B1(n1977), .B2(n17931), .ZN(
        n3035) );
  OAI22_X1 U1754 ( .A1(n18627), .A2(n18951), .B1(n1977), .B2(n17932), .ZN(
        n3036) );
  OAI22_X1 U1755 ( .A1(n18627), .A2(n18954), .B1(n18623), .B2(n17933), .ZN(
        n3037) );
  OAI22_X1 U1756 ( .A1(n18627), .A2(n18957), .B1(n18623), .B2(n17934), .ZN(
        n3038) );
  OAI22_X1 U1757 ( .A1(n18626), .A2(n18960), .B1(n18623), .B2(n17935), .ZN(
        n3039) );
  OAI22_X1 U1758 ( .A1(n1419), .A2(n18635), .B1(n18634), .B2(n17386), .ZN(
        n3051) );
  OAI22_X1 U1759 ( .A1(n1694), .A2(n18635), .B1(n18634), .B2(n17387), .ZN(
        n3052) );
  OAI22_X1 U1760 ( .A1(n18642), .A2(n18906), .B1(n18634), .B2(n17388), .ZN(
        n3053) );
  OAI22_X1 U1761 ( .A1(n18642), .A2(n18909), .B1(n18634), .B2(n17389), .ZN(
        n3054) );
  OAI22_X1 U1762 ( .A1(n18641), .A2(n18912), .B1(n18634), .B2(n17390), .ZN(
        n3055) );
  OAI22_X1 U1763 ( .A1(n18641), .A2(n18915), .B1(n18634), .B2(n17367), .ZN(
        n3056) );
  OAI22_X1 U1764 ( .A1(n18641), .A2(n18918), .B1(n18634), .B2(n17368), .ZN(
        n3057) );
  OAI22_X1 U1765 ( .A1(n18641), .A2(n18921), .B1(n18634), .B2(n17369), .ZN(
        n3058) );
  OAI22_X1 U1766 ( .A1(n18640), .A2(n18924), .B1(n18634), .B2(n17370), .ZN(
        n3059) );
  OAI22_X1 U1767 ( .A1(n18640), .A2(n18927), .B1(n1942), .B2(n17371), .ZN(
        n3060) );
  OAI22_X1 U1768 ( .A1(n18640), .A2(n18930), .B1(n1942), .B2(n17372), .ZN(
        n3061) );
  OAI22_X1 U1769 ( .A1(n18640), .A2(n18933), .B1(n1942), .B2(n17373), .ZN(
        n3062) );
  OAI22_X1 U1770 ( .A1(n18639), .A2(n18936), .B1(n1942), .B2(n17374), .ZN(
        n3063) );
  OAI22_X1 U1771 ( .A1(n18639), .A2(n18939), .B1(n1942), .B2(n17375), .ZN(
        n3064) );
  OAI22_X1 U1772 ( .A1(n18639), .A2(n18942), .B1(n1942), .B2(n17376), .ZN(
        n3065) );
  OAI22_X1 U1773 ( .A1(n18638), .A2(n18945), .B1(n1942), .B2(n17377), .ZN(
        n3066) );
  OAI22_X1 U1774 ( .A1(n18638), .A2(n18948), .B1(n1942), .B2(n17378), .ZN(
        n3067) );
  OAI22_X1 U1775 ( .A1(n18638), .A2(n18951), .B1(n1942), .B2(n17379), .ZN(
        n3068) );
  OAI22_X1 U1776 ( .A1(n18638), .A2(n18954), .B1(n18634), .B2(n17380), .ZN(
        n3069) );
  OAI22_X1 U1777 ( .A1(n18637), .A2(n18957), .B1(n18634), .B2(n17381), .ZN(
        n3070) );
  OAI22_X1 U1778 ( .A1(n18637), .A2(n18960), .B1(n18634), .B2(n17382), .ZN(
        n3071) );
  OAI22_X1 U1779 ( .A1(n1209), .A2(n18660), .B1(n18659), .B2(n17785), .ZN(
        n3113) );
  OAI22_X1 U1780 ( .A1(n1282), .A2(n18660), .B1(n18659), .B2(n17786), .ZN(
        n3114) );
  OAI22_X1 U1781 ( .A1(n1694), .A2(n18660), .B1(n18659), .B2(n17787), .ZN(
        n3116) );
  OAI22_X1 U1782 ( .A1(n18667), .A2(n18905), .B1(n18659), .B2(n17788), .ZN(
        n3117) );
  OAI22_X1 U1783 ( .A1(n18667), .A2(n18908), .B1(n18659), .B2(n17789), .ZN(
        n3118) );
  OAI22_X1 U1784 ( .A1(n18667), .A2(n18911), .B1(n18659), .B2(n17790), .ZN(
        n3119) );
  OAI22_X1 U1785 ( .A1(n18666), .A2(n18914), .B1(n18659), .B2(n17791), .ZN(
        n3120) );
  OAI22_X1 U1786 ( .A1(n18666), .A2(n18917), .B1(n18659), .B2(n17792), .ZN(
        n3121) );
  OAI22_X1 U1787 ( .A1(n18666), .A2(n18920), .B1(n18659), .B2(n17793), .ZN(
        n3122) );
  OAI22_X1 U1788 ( .A1(n18666), .A2(n18923), .B1(n18659), .B2(n17794), .ZN(
        n3123) );
  OAI22_X1 U1789 ( .A1(n18665), .A2(n18926), .B1(n1874), .B2(n17795), .ZN(
        n3124) );
  OAI22_X1 U1790 ( .A1(n18665), .A2(n18929), .B1(n1874), .B2(n17796), .ZN(
        n3125) );
  OAI22_X1 U1791 ( .A1(n18665), .A2(n18932), .B1(n1874), .B2(n17797), .ZN(
        n3126) );
  OAI22_X1 U1792 ( .A1(n18665), .A2(n18935), .B1(n1874), .B2(n17798), .ZN(
        n3127) );
  OAI22_X1 U1793 ( .A1(n18664), .A2(n18938), .B1(n1874), .B2(n17799), .ZN(
        n3128) );
  OAI22_X1 U1794 ( .A1(n18664), .A2(n18941), .B1(n1874), .B2(n17800), .ZN(
        n3129) );
  OAI22_X1 U1795 ( .A1(n18664), .A2(n18944), .B1(n1874), .B2(n17801), .ZN(
        n3130) );
  OAI22_X1 U1796 ( .A1(n18663), .A2(n18947), .B1(n1874), .B2(n17802), .ZN(
        n3131) );
  OAI22_X1 U1797 ( .A1(n18663), .A2(n18950), .B1(n1874), .B2(n17803), .ZN(
        n3132) );
  OAI22_X1 U1798 ( .A1(n18663), .A2(n18953), .B1(n18659), .B2(n17804), .ZN(
        n3133) );
  OAI22_X1 U1799 ( .A1(n18663), .A2(n18956), .B1(n18659), .B2(n17805), .ZN(
        n3134) );
  OAI22_X1 U1800 ( .A1(n18662), .A2(n18959), .B1(n18659), .B2(n17806), .ZN(
        n3135) );
  OAI22_X1 U1801 ( .A1(n1174), .A2(n18671), .B1(n18670), .B2(n17669), .ZN(
        n3144) );
  OAI22_X1 U1802 ( .A1(n1282), .A2(n18671), .B1(n18670), .B2(n17671), .ZN(
        n3146) );
  OAI22_X1 U1803 ( .A1(n1694), .A2(n18671), .B1(n18670), .B2(n17673), .ZN(
        n3148) );
  OAI22_X1 U1804 ( .A1(n18678), .A2(n18905), .B1(n18670), .B2(n17674), .ZN(
        n3149) );
  OAI22_X1 U1805 ( .A1(n18678), .A2(n18908), .B1(n18670), .B2(n17675), .ZN(
        n3150) );
  OAI22_X1 U1806 ( .A1(n18678), .A2(n18911), .B1(n18670), .B2(n17676), .ZN(
        n3151) );
  OAI22_X1 U1807 ( .A1(n18677), .A2(n18914), .B1(n18670), .B2(n17622), .ZN(
        n3152) );
  OAI22_X1 U1808 ( .A1(n18677), .A2(n18917), .B1(n18670), .B2(n17623), .ZN(
        n3153) );
  OAI22_X1 U1809 ( .A1(n18677), .A2(n18920), .B1(n18670), .B2(n17624), .ZN(
        n3154) );
  OAI22_X1 U1810 ( .A1(n18677), .A2(n18923), .B1(n18670), .B2(n17625), .ZN(
        n3155) );
  OAI22_X1 U1811 ( .A1(n18676), .A2(n18926), .B1(n1840), .B2(n17626), .ZN(
        n3156) );
  OAI22_X1 U1812 ( .A1(n18676), .A2(n18929), .B1(n1840), .B2(n17627), .ZN(
        n3157) );
  OAI22_X1 U1813 ( .A1(n18676), .A2(n18932), .B1(n1840), .B2(n17628), .ZN(
        n3158) );
  OAI22_X1 U1814 ( .A1(n18676), .A2(n18935), .B1(n1840), .B2(n17629), .ZN(
        n3159) );
  OAI22_X1 U1815 ( .A1(n18675), .A2(n18938), .B1(n1840), .B2(n17630), .ZN(
        n3160) );
  OAI22_X1 U1816 ( .A1(n18675), .A2(n18941), .B1(n1840), .B2(n17631), .ZN(
        n3161) );
  OAI22_X1 U1817 ( .A1(n18675), .A2(n18944), .B1(n1840), .B2(n17632), .ZN(
        n3162) );
  OAI22_X1 U1818 ( .A1(n18674), .A2(n18947), .B1(n1840), .B2(n17633), .ZN(
        n3163) );
  OAI22_X1 U1819 ( .A1(n18674), .A2(n18950), .B1(n1840), .B2(n17634), .ZN(
        n3164) );
  OAI22_X1 U1820 ( .A1(n18674), .A2(n18953), .B1(n18670), .B2(n17635), .ZN(
        n3165) );
  OAI22_X1 U1821 ( .A1(n18674), .A2(n18956), .B1(n18670), .B2(n17636), .ZN(
        n3166) );
  OAI22_X1 U1822 ( .A1(n18673), .A2(n18959), .B1(n18670), .B2(n17637), .ZN(
        n3167) );
  OAI22_X1 U1823 ( .A1(n1174), .A2(n18693), .B1(n18692), .B2(n18138), .ZN(
        n3208) );
  OAI22_X1 U1824 ( .A1(n1209), .A2(n18693), .B1(n18692), .B2(n18139), .ZN(
        n3209) );
  OAI22_X1 U1825 ( .A1(n1694), .A2(n18693), .B1(n18692), .B2(n18140), .ZN(
        n3212) );
  OAI22_X1 U1826 ( .A1(n18700), .A2(n18905), .B1(n18692), .B2(n18141), .ZN(
        n3213) );
  OAI22_X1 U1827 ( .A1(n18700), .A2(n18908), .B1(n18692), .B2(n18142), .ZN(
        n3214) );
  OAI22_X1 U1828 ( .A1(n18700), .A2(n18911), .B1(n18692), .B2(n18143), .ZN(
        n3215) );
  OAI22_X1 U1829 ( .A1(n18699), .A2(n18914), .B1(n18692), .B2(n18144), .ZN(
        n3216) );
  OAI22_X1 U1830 ( .A1(n18699), .A2(n18917), .B1(n18692), .B2(n18145), .ZN(
        n3217) );
  OAI22_X1 U1831 ( .A1(n18699), .A2(n18920), .B1(n18692), .B2(n18146), .ZN(
        n3218) );
  OAI22_X1 U1832 ( .A1(n18699), .A2(n18923), .B1(n18692), .B2(n18147), .ZN(
        n3219) );
  OAI22_X1 U1833 ( .A1(n18698), .A2(n18926), .B1(n1770), .B2(n18148), .ZN(
        n3220) );
  OAI22_X1 U1834 ( .A1(n18698), .A2(n18929), .B1(n1770), .B2(n18149), .ZN(
        n3221) );
  OAI22_X1 U1835 ( .A1(n18698), .A2(n18932), .B1(n1770), .B2(n18150), .ZN(
        n3222) );
  OAI22_X1 U1836 ( .A1(n18698), .A2(n18935), .B1(n1770), .B2(n18151), .ZN(
        n3223) );
  OAI22_X1 U1837 ( .A1(n18697), .A2(n18938), .B1(n1770), .B2(n18152), .ZN(
        n3224) );
  OAI22_X1 U1838 ( .A1(n18697), .A2(n18941), .B1(n1770), .B2(n18153), .ZN(
        n3225) );
  OAI22_X1 U1839 ( .A1(n18697), .A2(n18944), .B1(n1770), .B2(n18154), .ZN(
        n3226) );
  OAI22_X1 U1840 ( .A1(n18696), .A2(n18947), .B1(n1770), .B2(n18155), .ZN(
        n3227) );
  OAI22_X1 U1841 ( .A1(n18696), .A2(n18950), .B1(n1770), .B2(n18156), .ZN(
        n3228) );
  OAI22_X1 U1842 ( .A1(n18696), .A2(n18953), .B1(n18692), .B2(n18157), .ZN(
        n3229) );
  OAI22_X1 U1843 ( .A1(n18696), .A2(n18956), .B1(n18692), .B2(n18158), .ZN(
        n3230) );
  OAI22_X1 U1844 ( .A1(n18695), .A2(n18959), .B1(n18692), .B2(n18159), .ZN(
        n3231) );
  OAI22_X1 U1845 ( .A1(n1209), .A2(n18704), .B1(n18703), .B2(n17883), .ZN(
        n3241) );
  OAI22_X1 U1846 ( .A1(n1694), .A2(n18704), .B1(n18703), .B2(n17884), .ZN(
        n3244) );
  OAI22_X1 U1847 ( .A1(n18711), .A2(n18905), .B1(n18703), .B2(n17885), .ZN(
        n3245) );
  OAI22_X1 U1848 ( .A1(n18711), .A2(n18908), .B1(n18703), .B2(n17886), .ZN(
        n3246) );
  OAI22_X1 U1849 ( .A1(n18710), .A2(n18911), .B1(n18703), .B2(n17887), .ZN(
        n3247) );
  OAI22_X1 U1850 ( .A1(n18710), .A2(n18914), .B1(n18703), .B2(n17888), .ZN(
        n3248) );
  OAI22_X1 U1851 ( .A1(n18710), .A2(n18917), .B1(n18703), .B2(n17889), .ZN(
        n3249) );
  OAI22_X1 U1852 ( .A1(n18710), .A2(n18920), .B1(n18703), .B2(n17890), .ZN(
        n3250) );
  OAI22_X1 U1853 ( .A1(n18709), .A2(n18923), .B1(n18703), .B2(n17891), .ZN(
        n3251) );
  OAI22_X1 U1854 ( .A1(n18709), .A2(n18926), .B1(n1736), .B2(n17892), .ZN(
        n3252) );
  OAI22_X1 U1855 ( .A1(n18709), .A2(n18929), .B1(n1736), .B2(n17893), .ZN(
        n3253) );
  OAI22_X1 U1856 ( .A1(n18709), .A2(n18932), .B1(n1736), .B2(n17894), .ZN(
        n3254) );
  OAI22_X1 U1857 ( .A1(n18708), .A2(n18935), .B1(n1736), .B2(n17895), .ZN(
        n3255) );
  OAI22_X1 U1858 ( .A1(n18708), .A2(n18938), .B1(n1736), .B2(n17896), .ZN(
        n3256) );
  OAI22_X1 U1859 ( .A1(n18708), .A2(n18941), .B1(n1736), .B2(n17897), .ZN(
        n3257) );
  OAI22_X1 U1860 ( .A1(n18707), .A2(n18944), .B1(n1736), .B2(n17898), .ZN(
        n3258) );
  OAI22_X1 U1861 ( .A1(n18707), .A2(n18947), .B1(n1736), .B2(n17899), .ZN(
        n3259) );
  OAI22_X1 U1862 ( .A1(n18707), .A2(n18950), .B1(n1736), .B2(n17900), .ZN(
        n3260) );
  OAI22_X1 U1863 ( .A1(n18707), .A2(n18953), .B1(n18703), .B2(n17901), .ZN(
        n3261) );
  OAI22_X1 U1864 ( .A1(n18706), .A2(n18956), .B1(n18703), .B2(n17902), .ZN(
        n3262) );
  OAI22_X1 U1865 ( .A1(n18706), .A2(n18959), .B1(n18703), .B2(n17903), .ZN(
        n3263) );
  OAI22_X1 U1866 ( .A1(n1174), .A2(n18715), .B1(n18714), .B2(n17754), .ZN(
        n3272) );
  OAI22_X1 U1867 ( .A1(n1694), .A2(n18715), .B1(n18714), .B2(n17755), .ZN(
        n3276) );
  OAI22_X1 U1868 ( .A1(n18722), .A2(n18905), .B1(n18714), .B2(n17756), .ZN(
        n3277) );
  OAI22_X1 U1869 ( .A1(n18722), .A2(n18908), .B1(n18714), .B2(n17757), .ZN(
        n3278) );
  OAI22_X1 U1870 ( .A1(n18721), .A2(n18911), .B1(n18714), .B2(n17758), .ZN(
        n3279) );
  OAI22_X1 U1871 ( .A1(n18721), .A2(n18914), .B1(n18714), .B2(n17759), .ZN(
        n3280) );
  OAI22_X1 U1872 ( .A1(n18721), .A2(n18917), .B1(n18714), .B2(n17760), .ZN(
        n3281) );
  OAI22_X1 U1873 ( .A1(n18721), .A2(n18920), .B1(n18714), .B2(n17761), .ZN(
        n3282) );
  OAI22_X1 U1874 ( .A1(n18720), .A2(n18923), .B1(n18714), .B2(n17762), .ZN(
        n3283) );
  OAI22_X1 U1875 ( .A1(n18720), .A2(n18926), .B1(n1702), .B2(n17763), .ZN(
        n3284) );
  OAI22_X1 U1876 ( .A1(n18720), .A2(n18929), .B1(n1702), .B2(n17764), .ZN(
        n3285) );
  OAI22_X1 U1877 ( .A1(n18720), .A2(n18932), .B1(n1702), .B2(n17765), .ZN(
        n3286) );
  OAI22_X1 U1878 ( .A1(n18719), .A2(n18935), .B1(n1702), .B2(n17766), .ZN(
        n3287) );
  OAI22_X1 U1879 ( .A1(n18719), .A2(n18938), .B1(n1702), .B2(n17767), .ZN(
        n3288) );
  OAI22_X1 U1880 ( .A1(n18719), .A2(n18941), .B1(n1702), .B2(n17768), .ZN(
        n3289) );
  OAI22_X1 U1881 ( .A1(n18718), .A2(n18944), .B1(n1702), .B2(n17769), .ZN(
        n3290) );
  OAI22_X1 U1882 ( .A1(n18718), .A2(n18947), .B1(n1702), .B2(n17770), .ZN(
        n3291) );
  OAI22_X1 U1883 ( .A1(n18718), .A2(n18950), .B1(n1702), .B2(n17771), .ZN(
        n3292) );
  OAI22_X1 U1884 ( .A1(n18718), .A2(n18953), .B1(n18714), .B2(n17772), .ZN(
        n3293) );
  OAI22_X1 U1885 ( .A1(n18717), .A2(n18956), .B1(n18714), .B2(n17773), .ZN(
        n3294) );
  OAI22_X1 U1886 ( .A1(n18717), .A2(n18959), .B1(n18714), .B2(n17774), .ZN(
        n3295) );
  OAI22_X1 U1887 ( .A1(n1694), .A2(n18726), .B1(n18725), .B2(n18086), .ZN(
        n3308) );
  OAI22_X1 U1888 ( .A1(n18733), .A2(n18905), .B1(n18725), .B2(n18087), .ZN(
        n3309) );
  OAI22_X1 U1889 ( .A1(n18732), .A2(n18908), .B1(n18725), .B2(n18088), .ZN(
        n3310) );
  OAI22_X1 U1890 ( .A1(n18732), .A2(n18911), .B1(n18725), .B2(n18089), .ZN(
        n3311) );
  OAI22_X1 U1891 ( .A1(n18732), .A2(n18914), .B1(n18725), .B2(n18090), .ZN(
        n3312) );
  OAI22_X1 U1892 ( .A1(n18732), .A2(n18917), .B1(n18725), .B2(n18091), .ZN(
        n3313) );
  OAI22_X1 U1893 ( .A1(n18731), .A2(n18920), .B1(n18725), .B2(n18092), .ZN(
        n3314) );
  OAI22_X1 U1894 ( .A1(n18731), .A2(n18923), .B1(n18725), .B2(n18093), .ZN(
        n3315) );
  OAI22_X1 U1895 ( .A1(n18731), .A2(n18926), .B1(n1666), .B2(n18094), .ZN(
        n3316) );
  OAI22_X1 U1896 ( .A1(n18731), .A2(n18929), .B1(n1666), .B2(n18095), .ZN(
        n3317) );
  OAI22_X1 U1897 ( .A1(n18730), .A2(n18932), .B1(n1666), .B2(n18096), .ZN(
        n3318) );
  OAI22_X1 U1898 ( .A1(n18730), .A2(n18935), .B1(n1666), .B2(n18097), .ZN(
        n3319) );
  OAI22_X1 U1899 ( .A1(n18730), .A2(n18938), .B1(n1666), .B2(n18098), .ZN(
        n3320) );
  OAI22_X1 U1900 ( .A1(n18729), .A2(n18941), .B1(n1666), .B2(n18099), .ZN(
        n3321) );
  OAI22_X1 U1901 ( .A1(n18729), .A2(n18944), .B1(n1666), .B2(n18100), .ZN(
        n3322) );
  OAI22_X1 U1902 ( .A1(n18729), .A2(n18947), .B1(n1666), .B2(n18101), .ZN(
        n3323) );
  OAI22_X1 U1903 ( .A1(n18729), .A2(n18950), .B1(n1666), .B2(n18102), .ZN(
        n3324) );
  OAI22_X1 U1904 ( .A1(n18728), .A2(n18953), .B1(n18725), .B2(n18103), .ZN(
        n3325) );
  OAI22_X1 U1905 ( .A1(n18728), .A2(n18956), .B1(n18725), .B2(n18104), .ZN(
        n3326) );
  OAI22_X1 U1906 ( .A1(n18728), .A2(n18959), .B1(n18725), .B2(n18105), .ZN(
        n3327) );
  OAI22_X1 U1907 ( .A1(n1209), .A2(n18751), .B1(n18750), .B2(n17849), .ZN(
        n3369) );
  OAI22_X1 U1908 ( .A1(n1282), .A2(n18751), .B1(n18750), .B2(n17850), .ZN(
        n3370) );
  OAI22_X1 U1909 ( .A1(n1419), .A2(n18751), .B1(n18750), .B2(n17851), .ZN(
        n3371) );
  OAI22_X1 U1910 ( .A1(n18758), .A2(n18905), .B1(n18750), .B2(n17853), .ZN(
        n3373) );
  OAI22_X1 U1911 ( .A1(n18758), .A2(n18908), .B1(n18750), .B2(n17854), .ZN(
        n3374) );
  OAI22_X1 U1912 ( .A1(n18758), .A2(n18911), .B1(n18750), .B2(n17855), .ZN(
        n3375) );
  OAI22_X1 U1913 ( .A1(n18757), .A2(n18914), .B1(n18750), .B2(n17856), .ZN(
        n3376) );
  OAI22_X1 U1914 ( .A1(n18757), .A2(n18917), .B1(n18750), .B2(n17857), .ZN(
        n3377) );
  OAI22_X1 U1915 ( .A1(n18757), .A2(n18920), .B1(n18750), .B2(n17858), .ZN(
        n3378) );
  OAI22_X1 U1916 ( .A1(n18757), .A2(n18923), .B1(n18750), .B2(n17859), .ZN(
        n3379) );
  OAI22_X1 U1917 ( .A1(n18756), .A2(n18926), .B1(n1597), .B2(n17860), .ZN(
        n3380) );
  OAI22_X1 U1918 ( .A1(n18756), .A2(n18929), .B1(n1597), .B2(n17861), .ZN(
        n3381) );
  OAI22_X1 U1919 ( .A1(n18756), .A2(n18932), .B1(n1597), .B2(n17862), .ZN(
        n3382) );
  OAI22_X1 U1920 ( .A1(n18756), .A2(n18935), .B1(n1597), .B2(n17863), .ZN(
        n3383) );
  OAI22_X1 U1921 ( .A1(n18755), .A2(n18938), .B1(n1597), .B2(n17864), .ZN(
        n3384) );
  OAI22_X1 U1922 ( .A1(n18755), .A2(n18941), .B1(n1597), .B2(n17865), .ZN(
        n3385) );
  OAI22_X1 U1923 ( .A1(n18755), .A2(n18944), .B1(n1597), .B2(n17866), .ZN(
        n3386) );
  OAI22_X1 U1924 ( .A1(n18754), .A2(n18947), .B1(n1597), .B2(n17867), .ZN(
        n3387) );
  OAI22_X1 U1925 ( .A1(n18754), .A2(n18950), .B1(n18750), .B2(n17868), .ZN(
        n3388) );
  OAI22_X1 U1926 ( .A1(n18754), .A2(n18953), .B1(n18750), .B2(n17869), .ZN(
        n3389) );
  OAI22_X1 U1927 ( .A1(n18754), .A2(n18956), .B1(n18750), .B2(n17870), .ZN(
        n3390) );
  OAI22_X1 U1928 ( .A1(n18753), .A2(n18959), .B1(n18750), .B2(n17871), .ZN(
        n3391) );
  OAI22_X1 U1929 ( .A1(n1174), .A2(n18762), .B1(n18761), .B2(n18170), .ZN(
        n3400) );
  OAI22_X1 U1930 ( .A1(n1282), .A2(n18762), .B1(n18761), .B2(n18171), .ZN(
        n3402) );
  OAI22_X1 U1931 ( .A1(n1419), .A2(n18762), .B1(n18761), .B2(n18172), .ZN(
        n3403) );
  OAI22_X1 U1932 ( .A1(n18769), .A2(n18905), .B1(n18761), .B2(n18173), .ZN(
        n3405) );
  OAI22_X1 U1933 ( .A1(n18769), .A2(n18908), .B1(n18761), .B2(n18174), .ZN(
        n3406) );
  OAI22_X1 U1934 ( .A1(n18769), .A2(n18911), .B1(n18761), .B2(n18175), .ZN(
        n3407) );
  OAI22_X1 U1935 ( .A1(n18768), .A2(n18914), .B1(n18761), .B2(n18176), .ZN(
        n3408) );
  OAI22_X1 U1936 ( .A1(n18768), .A2(n18917), .B1(n18761), .B2(n18177), .ZN(
        n3409) );
  OAI22_X1 U1937 ( .A1(n18768), .A2(n18920), .B1(n18761), .B2(n18178), .ZN(
        n3410) );
  OAI22_X1 U1938 ( .A1(n18768), .A2(n18923), .B1(n18761), .B2(n18179), .ZN(
        n3411) );
  OAI22_X1 U1939 ( .A1(n18767), .A2(n18926), .B1(n1563), .B2(n18180), .ZN(
        n3412) );
  OAI22_X1 U1940 ( .A1(n18767), .A2(n18929), .B1(n1563), .B2(n18181), .ZN(
        n3413) );
  OAI22_X1 U1941 ( .A1(n18767), .A2(n18932), .B1(n1563), .B2(n18182), .ZN(
        n3414) );
  OAI22_X1 U1942 ( .A1(n18767), .A2(n18935), .B1(n1563), .B2(n18183), .ZN(
        n3415) );
  OAI22_X1 U1943 ( .A1(n18766), .A2(n18938), .B1(n1563), .B2(n18184), .ZN(
        n3416) );
  OAI22_X1 U1944 ( .A1(n18766), .A2(n18941), .B1(n1563), .B2(n18185), .ZN(
        n3417) );
  OAI22_X1 U1945 ( .A1(n18766), .A2(n18944), .B1(n1563), .B2(n18186), .ZN(
        n3418) );
  OAI22_X1 U1946 ( .A1(n18765), .A2(n18947), .B1(n1563), .B2(n18187), .ZN(
        n3419) );
  OAI22_X1 U1947 ( .A1(n18765), .A2(n18950), .B1(n18761), .B2(n18188), .ZN(
        n3420) );
  OAI22_X1 U1948 ( .A1(n18765), .A2(n18953), .B1(n18761), .B2(n18189), .ZN(
        n3421) );
  OAI22_X1 U1949 ( .A1(n18765), .A2(n18956), .B1(n18761), .B2(n18190), .ZN(
        n3422) );
  OAI22_X1 U1950 ( .A1(n18764), .A2(n18959), .B1(n18761), .B2(n18191), .ZN(
        n3423) );
  OAI22_X1 U1951 ( .A1(n1282), .A2(n18773), .B1(n18772), .B2(n18022), .ZN(
        n3434) );
  OAI22_X1 U1952 ( .A1(n1419), .A2(n18773), .B1(n18772), .B2(n18023), .ZN(
        n3435) );
  OAI22_X1 U1953 ( .A1(n18780), .A2(n18905), .B1(n18772), .B2(n18024), .ZN(
        n3437) );
  OAI22_X1 U1954 ( .A1(n18780), .A2(n18908), .B1(n18772), .B2(n18025), .ZN(
        n3438) );
  OAI22_X1 U1955 ( .A1(n18779), .A2(n18911), .B1(n18772), .B2(n18026), .ZN(
        n3439) );
  OAI22_X1 U1956 ( .A1(n18779), .A2(n18914), .B1(n18772), .B2(n18027), .ZN(
        n3440) );
  OAI22_X1 U1957 ( .A1(n18779), .A2(n18917), .B1(n18772), .B2(n18028), .ZN(
        n3441) );
  OAI22_X1 U1958 ( .A1(n18779), .A2(n18920), .B1(n18772), .B2(n18029), .ZN(
        n3442) );
  OAI22_X1 U1959 ( .A1(n18778), .A2(n18923), .B1(n18772), .B2(n18030), .ZN(
        n3443) );
  OAI22_X1 U1960 ( .A1(n18778), .A2(n18926), .B1(n1528), .B2(n18031), .ZN(
        n3444) );
  OAI22_X1 U1961 ( .A1(n18778), .A2(n18929), .B1(n1528), .B2(n18032), .ZN(
        n3445) );
  OAI22_X1 U1962 ( .A1(n18778), .A2(n18932), .B1(n1528), .B2(n18033), .ZN(
        n3446) );
  OAI22_X1 U1963 ( .A1(n18777), .A2(n18935), .B1(n1528), .B2(n18034), .ZN(
        n3447) );
  OAI22_X1 U1964 ( .A1(n18777), .A2(n18938), .B1(n1528), .B2(n18035), .ZN(
        n3448) );
  OAI22_X1 U1965 ( .A1(n18777), .A2(n18941), .B1(n1528), .B2(n18036), .ZN(
        n3449) );
  OAI22_X1 U1966 ( .A1(n18776), .A2(n18944), .B1(n1528), .B2(n18037), .ZN(
        n3450) );
  OAI22_X1 U1967 ( .A1(n18776), .A2(n18947), .B1(n1528), .B2(n18038), .ZN(
        n3451) );
  OAI22_X1 U1968 ( .A1(n18776), .A2(n18950), .B1(n18772), .B2(n18039), .ZN(
        n3452) );
  OAI22_X1 U1969 ( .A1(n18776), .A2(n18953), .B1(n18772), .B2(n18040), .ZN(
        n3453) );
  OAI22_X1 U1970 ( .A1(n18775), .A2(n18956), .B1(n18772), .B2(n18041), .ZN(
        n3454) );
  OAI22_X1 U1971 ( .A1(n18775), .A2(n18959), .B1(n18772), .B2(n18042), .ZN(
        n3455) );
  OAI22_X1 U1972 ( .A1(n1174), .A2(n18784), .B1(n18783), .B2(n18106), .ZN(
        n3464) );
  OAI22_X1 U1973 ( .A1(n1209), .A2(n18784), .B1(n18783), .B2(n18107), .ZN(
        n3465) );
  OAI22_X1 U1974 ( .A1(n1419), .A2(n18784), .B1(n18783), .B2(n18108), .ZN(
        n3467) );
  OAI22_X1 U1975 ( .A1(n18791), .A2(n18904), .B1(n18783), .B2(n18109), .ZN(
        n3469) );
  OAI22_X1 U1976 ( .A1(n18791), .A2(n18907), .B1(n18783), .B2(n18110), .ZN(
        n3470) );
  OAI22_X1 U1977 ( .A1(n18791), .A2(n18910), .B1(n18783), .B2(n18111), .ZN(
        n3471) );
  OAI22_X1 U1978 ( .A1(n18790), .A2(n18913), .B1(n18783), .B2(n18112), .ZN(
        n3472) );
  OAI22_X1 U1979 ( .A1(n18790), .A2(n18916), .B1(n18783), .B2(n18113), .ZN(
        n3473) );
  OAI22_X1 U1980 ( .A1(n18790), .A2(n18919), .B1(n18783), .B2(n18114), .ZN(
        n3474) );
  OAI22_X1 U1981 ( .A1(n18790), .A2(n18922), .B1(n18783), .B2(n18115), .ZN(
        n3475) );
  OAI22_X1 U1982 ( .A1(n18789), .A2(n18925), .B1(n1494), .B2(n18116), .ZN(
        n3476) );
  OAI22_X1 U1983 ( .A1(n18789), .A2(n18928), .B1(n1494), .B2(n18117), .ZN(
        n3477) );
  OAI22_X1 U1984 ( .A1(n18789), .A2(n18931), .B1(n1494), .B2(n18118), .ZN(
        n3478) );
  OAI22_X1 U1985 ( .A1(n18789), .A2(n18934), .B1(n1494), .B2(n18119), .ZN(
        n3479) );
  OAI22_X1 U1986 ( .A1(n18788), .A2(n18937), .B1(n1494), .B2(n18120), .ZN(
        n3480) );
  OAI22_X1 U1987 ( .A1(n18788), .A2(n18940), .B1(n1494), .B2(n18121), .ZN(
        n3481) );
  OAI22_X1 U1988 ( .A1(n18788), .A2(n18943), .B1(n1494), .B2(n18122), .ZN(
        n3482) );
  OAI22_X1 U1989 ( .A1(n18787), .A2(n18946), .B1(n1494), .B2(n18123), .ZN(
        n3483) );
  OAI22_X1 U1990 ( .A1(n18787), .A2(n18949), .B1(n18783), .B2(n18124), .ZN(
        n3484) );
  OAI22_X1 U1991 ( .A1(n18787), .A2(n18952), .B1(n18783), .B2(n18125), .ZN(
        n3485) );
  OAI22_X1 U1992 ( .A1(n18787), .A2(n18955), .B1(n18783), .B2(n18126), .ZN(
        n3486) );
  OAI22_X1 U1993 ( .A1(n18786), .A2(n18958), .B1(n18783), .B2(n18127), .ZN(
        n3487) );
  OAI22_X1 U1994 ( .A1(n1209), .A2(n18795), .B1(n18794), .B2(n17562), .ZN(
        n3497) );
  OAI22_X1 U1995 ( .A1(n1419), .A2(n18795), .B1(n18794), .B2(n17563), .ZN(
        n3499) );
  OAI22_X1 U1996 ( .A1(n18802), .A2(n18904), .B1(n18794), .B2(n17564), .ZN(
        n3501) );
  OAI22_X1 U1997 ( .A1(n18802), .A2(n18907), .B1(n18794), .B2(n17565), .ZN(
        n3502) );
  OAI22_X1 U1998 ( .A1(n18801), .A2(n18910), .B1(n18794), .B2(n17566), .ZN(
        n3503) );
  OAI22_X1 U1999 ( .A1(n18801), .A2(n18913), .B1(n18794), .B2(n17567), .ZN(
        n3504) );
  OAI22_X1 U2000 ( .A1(n18801), .A2(n18916), .B1(n18794), .B2(n17568), .ZN(
        n3505) );
  OAI22_X1 U2001 ( .A1(n18801), .A2(n18919), .B1(n18794), .B2(n17569), .ZN(
        n3506) );
  OAI22_X1 U2002 ( .A1(n18800), .A2(n18922), .B1(n18794), .B2(n17570), .ZN(
        n3507) );
  OAI22_X1 U2003 ( .A1(n18800), .A2(n18925), .B1(n1460), .B2(n17571), .ZN(
        n3508) );
  OAI22_X1 U2004 ( .A1(n18800), .A2(n18928), .B1(n1460), .B2(n17572), .ZN(
        n3509) );
  OAI22_X1 U2005 ( .A1(n18800), .A2(n18931), .B1(n1460), .B2(n17573), .ZN(
        n3510) );
  OAI22_X1 U2006 ( .A1(n18799), .A2(n18934), .B1(n1460), .B2(n17574), .ZN(
        n3511) );
  OAI22_X1 U2007 ( .A1(n18799), .A2(n18937), .B1(n1460), .B2(n17575), .ZN(
        n3512) );
  OAI22_X1 U2008 ( .A1(n18799), .A2(n18940), .B1(n1460), .B2(n17576), .ZN(
        n3513) );
  OAI22_X1 U2009 ( .A1(n18798), .A2(n18943), .B1(n1460), .B2(n17577), .ZN(
        n3514) );
  OAI22_X1 U2010 ( .A1(n18798), .A2(n18946), .B1(n1460), .B2(n17578), .ZN(
        n3515) );
  OAI22_X1 U2011 ( .A1(n18798), .A2(n18949), .B1(n18794), .B2(n17579), .ZN(
        n3516) );
  OAI22_X1 U2012 ( .A1(n18798), .A2(n18952), .B1(n18794), .B2(n17580), .ZN(
        n3517) );
  OAI22_X1 U2013 ( .A1(n18797), .A2(n18955), .B1(n18794), .B2(n17581), .ZN(
        n3518) );
  OAI22_X1 U2014 ( .A1(n18797), .A2(n18958), .B1(n18794), .B2(n17582), .ZN(
        n3519) );
  OAI22_X1 U2015 ( .A1(n1174), .A2(n18806), .B1(n18805), .B2(n17402), .ZN(
        n3528) );
  OAI22_X1 U2016 ( .A1(n1419), .A2(n18806), .B1(n18805), .B2(n17403), .ZN(
        n3531) );
  OAI22_X1 U2017 ( .A1(n18813), .A2(n18904), .B1(n18805), .B2(n17404), .ZN(
        n3533) );
  OAI22_X1 U2018 ( .A1(n18813), .A2(n18907), .B1(n18805), .B2(n17405), .ZN(
        n3534) );
  OAI22_X1 U2019 ( .A1(n18812), .A2(n18910), .B1(n18805), .B2(n17406), .ZN(
        n3535) );
  OAI22_X1 U2020 ( .A1(n18812), .A2(n18913), .B1(n18805), .B2(n17407), .ZN(
        n3536) );
  OAI22_X1 U2021 ( .A1(n18812), .A2(n18916), .B1(n18805), .B2(n17408), .ZN(
        n3537) );
  OAI22_X1 U2022 ( .A1(n18812), .A2(n18919), .B1(n18805), .B2(n17409), .ZN(
        n3538) );
  OAI22_X1 U2023 ( .A1(n18811), .A2(n18922), .B1(n18805), .B2(n17410), .ZN(
        n3539) );
  OAI22_X1 U2024 ( .A1(n18811), .A2(n18925), .B1(n1426), .B2(n17411), .ZN(
        n3540) );
  OAI22_X1 U2025 ( .A1(n18811), .A2(n18928), .B1(n1426), .B2(n17412), .ZN(
        n3541) );
  OAI22_X1 U2026 ( .A1(n18811), .A2(n18931), .B1(n1426), .B2(n17413), .ZN(
        n3542) );
  OAI22_X1 U2027 ( .A1(n18810), .A2(n18934), .B1(n1426), .B2(n17414), .ZN(
        n3543) );
  OAI22_X1 U2028 ( .A1(n18810), .A2(n18937), .B1(n1426), .B2(n17415), .ZN(
        n3544) );
  OAI22_X1 U2029 ( .A1(n18810), .A2(n18940), .B1(n1426), .B2(n17416), .ZN(
        n3545) );
  OAI22_X1 U2030 ( .A1(n18809), .A2(n18943), .B1(n1426), .B2(n17417), .ZN(
        n3546) );
  OAI22_X1 U2031 ( .A1(n18809), .A2(n18946), .B1(n1426), .B2(n17418), .ZN(
        n3547) );
  OAI22_X1 U2032 ( .A1(n18809), .A2(n18949), .B1(n18805), .B2(n17419), .ZN(
        n3548) );
  OAI22_X1 U2033 ( .A1(n18809), .A2(n18952), .B1(n18805), .B2(n17420), .ZN(
        n3549) );
  OAI22_X1 U2034 ( .A1(n18808), .A2(n18955), .B1(n18805), .B2(n17421), .ZN(
        n3550) );
  OAI22_X1 U2035 ( .A1(n18808), .A2(n18958), .B1(n18805), .B2(n17422), .ZN(
        n3551) );
  OAI22_X1 U2036 ( .A1(n1419), .A2(n18817), .B1(n18816), .B2(n17691), .ZN(
        n3563) );
  OAI22_X1 U2037 ( .A1(n18824), .A2(n18904), .B1(n18816), .B2(n17692), .ZN(
        n3565) );
  OAI22_X1 U2038 ( .A1(n18823), .A2(n18907), .B1(n18816), .B2(n17693), .ZN(
        n3566) );
  OAI22_X1 U2039 ( .A1(n18823), .A2(n18910), .B1(n18816), .B2(n17694), .ZN(
        n3567) );
  OAI22_X1 U2040 ( .A1(n18823), .A2(n18913), .B1(n18816), .B2(n17695), .ZN(
        n3568) );
  OAI22_X1 U2041 ( .A1(n18823), .A2(n18916), .B1(n18816), .B2(n17696), .ZN(
        n3569) );
  OAI22_X1 U2042 ( .A1(n18822), .A2(n18919), .B1(n18816), .B2(n17697), .ZN(
        n3570) );
  OAI22_X1 U2043 ( .A1(n18822), .A2(n18922), .B1(n18816), .B2(n17698), .ZN(
        n3571) );
  OAI22_X1 U2044 ( .A1(n18822), .A2(n18925), .B1(n1390), .B2(n17699), .ZN(
        n3572) );
  OAI22_X1 U2045 ( .A1(n18822), .A2(n18928), .B1(n1390), .B2(n17700), .ZN(
        n3573) );
  OAI22_X1 U2046 ( .A1(n18821), .A2(n18931), .B1(n1390), .B2(n17701), .ZN(
        n3574) );
  OAI22_X1 U2047 ( .A1(n18821), .A2(n18934), .B1(n1390), .B2(n17702), .ZN(
        n3575) );
  OAI22_X1 U2048 ( .A1(n18821), .A2(n18937), .B1(n1390), .B2(n17703), .ZN(
        n3576) );
  OAI22_X1 U2049 ( .A1(n18820), .A2(n18940), .B1(n1390), .B2(n17704), .ZN(
        n3577) );
  OAI22_X1 U2050 ( .A1(n18820), .A2(n18943), .B1(n1390), .B2(n17705), .ZN(
        n3578) );
  OAI22_X1 U2051 ( .A1(n18820), .A2(n18946), .B1(n1390), .B2(n17706), .ZN(
        n3579) );
  OAI22_X1 U2052 ( .A1(n18820), .A2(n18949), .B1(n18816), .B2(n17707), .ZN(
        n3580) );
  OAI22_X1 U2053 ( .A1(n18819), .A2(n18952), .B1(n18816), .B2(n17708), .ZN(
        n3581) );
  OAI22_X1 U2054 ( .A1(n18819), .A2(n18955), .B1(n18816), .B2(n17709), .ZN(
        n3582) );
  OAI22_X1 U2055 ( .A1(n18819), .A2(n18958), .B1(n18816), .B2(n17710), .ZN(
        n3583) );
  OAI22_X1 U2056 ( .A1(n1174), .A2(n18828), .B1(n18827), .B2(n17817), .ZN(
        n3592) );
  OAI22_X1 U2057 ( .A1(n1209), .A2(n18828), .B1(n18827), .B2(n17818), .ZN(
        n3593) );
  OAI22_X1 U2058 ( .A1(n1282), .A2(n18828), .B1(n18827), .B2(n17819), .ZN(
        n3594) );
  OAI22_X1 U2059 ( .A1(n18829), .A2(n18904), .B1(n18827), .B2(n17820), .ZN(
        n3597) );
  OAI22_X1 U2060 ( .A1(n18829), .A2(n18907), .B1(n18827), .B2(n17821), .ZN(
        n3598) );
  OAI22_X1 U2061 ( .A1(n18829), .A2(n18910), .B1(n18827), .B2(n17822), .ZN(
        n3599) );
  OAI22_X1 U2062 ( .A1(n18830), .A2(n18913), .B1(n18827), .B2(n17823), .ZN(
        n3600) );
  OAI22_X1 U2063 ( .A1(n18830), .A2(n18916), .B1(n18827), .B2(n17824), .ZN(
        n3601) );
  OAI22_X1 U2064 ( .A1(n18830), .A2(n18919), .B1(n18827), .B2(n17825), .ZN(
        n3602) );
  OAI22_X1 U2065 ( .A1(n18830), .A2(n18922), .B1(n18827), .B2(n17826), .ZN(
        n3603) );
  OAI22_X1 U2066 ( .A1(n18831), .A2(n18925), .B1(n1356), .B2(n17827), .ZN(
        n3604) );
  OAI22_X1 U2067 ( .A1(n18831), .A2(n18928), .B1(n1356), .B2(n17828), .ZN(
        n3605) );
  OAI22_X1 U2068 ( .A1(n18831), .A2(n18931), .B1(n1356), .B2(n17829), .ZN(
        n3606) );
  OAI22_X1 U2069 ( .A1(n18831), .A2(n18934), .B1(n1356), .B2(n17830), .ZN(
        n3607) );
  OAI22_X1 U2070 ( .A1(n18832), .A2(n18937), .B1(n1356), .B2(n17831), .ZN(
        n3608) );
  OAI22_X1 U2071 ( .A1(n18832), .A2(n18940), .B1(n1356), .B2(n17832), .ZN(
        n3609) );
  OAI22_X1 U2072 ( .A1(n18832), .A2(n18943), .B1(n1356), .B2(n17833), .ZN(
        n3610) );
  OAI22_X1 U2073 ( .A1(n18832), .A2(n18946), .B1(n1356), .B2(n17834), .ZN(
        n3611) );
  OAI22_X1 U2074 ( .A1(n18833), .A2(n18949), .B1(n18827), .B2(n17835), .ZN(
        n3612) );
  OAI22_X1 U2075 ( .A1(n18833), .A2(n18952), .B1(n18827), .B2(n17836), .ZN(
        n3613) );
  OAI22_X1 U2076 ( .A1(n18833), .A2(n18955), .B1(n18827), .B2(n17837), .ZN(
        n3614) );
  OAI22_X1 U2077 ( .A1(n18833), .A2(n18958), .B1(n18827), .B2(n17838), .ZN(
        n3615) );
  OAI22_X1 U2078 ( .A1(n1209), .A2(n18839), .B1(n18838), .B2(n17338), .ZN(
        n3625) );
  OAI22_X1 U2079 ( .A1(n1282), .A2(n18839), .B1(n18838), .B2(n17339), .ZN(
        n3626) );
  OAI22_X1 U2080 ( .A1(n18846), .A2(n18904), .B1(n18838), .B2(n17340), .ZN(
        n3629) );
  OAI22_X1 U2081 ( .A1(n18846), .A2(n18907), .B1(n18838), .B2(n17341), .ZN(
        n3630) );
  OAI22_X1 U2082 ( .A1(n18845), .A2(n18910), .B1(n18838), .B2(n17342), .ZN(
        n3631) );
  OAI22_X1 U2083 ( .A1(n18845), .A2(n18913), .B1(n18838), .B2(n17343), .ZN(
        n3632) );
  OAI22_X1 U2084 ( .A1(n18845), .A2(n18916), .B1(n18838), .B2(n17344), .ZN(
        n3633) );
  OAI22_X1 U2085 ( .A1(n18845), .A2(n18919), .B1(n18838), .B2(n17345), .ZN(
        n3634) );
  OAI22_X1 U2086 ( .A1(n18844), .A2(n18922), .B1(n18838), .B2(n17346), .ZN(
        n3635) );
  OAI22_X1 U2087 ( .A1(n18844), .A2(n18925), .B1(n1322), .B2(n17347), .ZN(
        n3636) );
  OAI22_X1 U2088 ( .A1(n18844), .A2(n18928), .B1(n1322), .B2(n17348), .ZN(
        n3637) );
  OAI22_X1 U2089 ( .A1(n18844), .A2(n18931), .B1(n1322), .B2(n17349), .ZN(
        n3638) );
  OAI22_X1 U2090 ( .A1(n18843), .A2(n18934), .B1(n1322), .B2(n17350), .ZN(
        n3639) );
  OAI22_X1 U2091 ( .A1(n18843), .A2(n18937), .B1(n1322), .B2(n17351), .ZN(
        n3640) );
  OAI22_X1 U2092 ( .A1(n18843), .A2(n18940), .B1(n1322), .B2(n17352), .ZN(
        n3641) );
  OAI22_X1 U2093 ( .A1(n18842), .A2(n18943), .B1(n1322), .B2(n17353), .ZN(
        n3642) );
  OAI22_X1 U2094 ( .A1(n18842), .A2(n18946), .B1(n1322), .B2(n17354), .ZN(
        n3643) );
  OAI22_X1 U2095 ( .A1(n18842), .A2(n18949), .B1(n18838), .B2(n17355), .ZN(
        n3644) );
  OAI22_X1 U2096 ( .A1(n18842), .A2(n18952), .B1(n18838), .B2(n17356), .ZN(
        n3645) );
  OAI22_X1 U2097 ( .A1(n18841), .A2(n18955), .B1(n18838), .B2(n17357), .ZN(
        n3646) );
  OAI22_X1 U2098 ( .A1(n18841), .A2(n18958), .B1(n18838), .B2(n17358), .ZN(
        n3647) );
  OAI22_X1 U2099 ( .A1(n1174), .A2(n18850), .B1(n18849), .B2(n18043), .ZN(
        n3656) );
  OAI22_X1 U2100 ( .A1(n1282), .A2(n18850), .B1(n18849), .B2(n18044), .ZN(
        n3658) );
  OAI22_X1 U2101 ( .A1(n18857), .A2(n18904), .B1(n18849), .B2(n18045), .ZN(
        n3661) );
  OAI22_X1 U2102 ( .A1(n18857), .A2(n18907), .B1(n18849), .B2(n18046), .ZN(
        n3662) );
  OAI22_X1 U2103 ( .A1(n18856), .A2(n18910), .B1(n18849), .B2(n18047), .ZN(
        n3663) );
  OAI22_X1 U2104 ( .A1(n18856), .A2(n18913), .B1(n18849), .B2(n18048), .ZN(
        n3664) );
  OAI22_X1 U2105 ( .A1(n18856), .A2(n18916), .B1(n18849), .B2(n18049), .ZN(
        n3665) );
  OAI22_X1 U2106 ( .A1(n18856), .A2(n18919), .B1(n18849), .B2(n18050), .ZN(
        n3666) );
  OAI22_X1 U2107 ( .A1(n18855), .A2(n18922), .B1(n18849), .B2(n18051), .ZN(
        n3667) );
  OAI22_X1 U2108 ( .A1(n18855), .A2(n18925), .B1(n1288), .B2(n18052), .ZN(
        n3668) );
  OAI22_X1 U2109 ( .A1(n18855), .A2(n18928), .B1(n1288), .B2(n18053), .ZN(
        n3669) );
  OAI22_X1 U2110 ( .A1(n18855), .A2(n18931), .B1(n1288), .B2(n18054), .ZN(
        n3670) );
  OAI22_X1 U2111 ( .A1(n18854), .A2(n18934), .B1(n1288), .B2(n18055), .ZN(
        n3671) );
  OAI22_X1 U2112 ( .A1(n18854), .A2(n18937), .B1(n1288), .B2(n18056), .ZN(
        n3672) );
  OAI22_X1 U2113 ( .A1(n18854), .A2(n18940), .B1(n1288), .B2(n18057), .ZN(
        n3673) );
  OAI22_X1 U2114 ( .A1(n18853), .A2(n18943), .B1(n1288), .B2(n18058), .ZN(
        n3674) );
  OAI22_X1 U2115 ( .A1(n18853), .A2(n18946), .B1(n1288), .B2(n18059), .ZN(
        n3675) );
  OAI22_X1 U2116 ( .A1(n18853), .A2(n18949), .B1(n18849), .B2(n18060), .ZN(
        n3676) );
  OAI22_X1 U2117 ( .A1(n18853), .A2(n18952), .B1(n18849), .B2(n18061), .ZN(
        n3677) );
  OAI22_X1 U2118 ( .A1(n18852), .A2(n18955), .B1(n18849), .B2(n18062), .ZN(
        n3678) );
  OAI22_X1 U2119 ( .A1(n18852), .A2(n18958), .B1(n18849), .B2(n18063), .ZN(
        n3679) );
  OAI22_X1 U2120 ( .A1(n1282), .A2(n18861), .B1(n18860), .B2(n18266), .ZN(
        n3690) );
  OAI22_X1 U2121 ( .A1(n18868), .A2(n18904), .B1(n18860), .B2(n18267), .ZN(
        n3693) );
  OAI22_X1 U2122 ( .A1(n18867), .A2(n18907), .B1(n18860), .B2(n18268), .ZN(
        n3694) );
  OAI22_X1 U2123 ( .A1(n18867), .A2(n18910), .B1(n18860), .B2(n18269), .ZN(
        n3695) );
  OAI22_X1 U2124 ( .A1(n18867), .A2(n18913), .B1(n18860), .B2(n18270), .ZN(
        n3696) );
  OAI22_X1 U2125 ( .A1(n18867), .A2(n18916), .B1(n18860), .B2(n18271), .ZN(
        n3697) );
  OAI22_X1 U2126 ( .A1(n18866), .A2(n18919), .B1(n18860), .B2(n18272), .ZN(
        n3698) );
  OAI22_X1 U2127 ( .A1(n18866), .A2(n18922), .B1(n18860), .B2(n18273), .ZN(
        n3699) );
  OAI22_X1 U2128 ( .A1(n18866), .A2(n18925), .B1(n1252), .B2(n18274), .ZN(
        n3700) );
  OAI22_X1 U2129 ( .A1(n18866), .A2(n18928), .B1(n1252), .B2(n18275), .ZN(
        n3701) );
  OAI22_X1 U2130 ( .A1(n18865), .A2(n18931), .B1(n1252), .B2(n18276), .ZN(
        n3702) );
  OAI22_X1 U2131 ( .A1(n18865), .A2(n18934), .B1(n1252), .B2(n18277), .ZN(
        n3703) );
  OAI22_X1 U2132 ( .A1(n18865), .A2(n18937), .B1(n1252), .B2(n18278), .ZN(
        n3704) );
  OAI22_X1 U2133 ( .A1(n18864), .A2(n18940), .B1(n1252), .B2(n18279), .ZN(
        n3705) );
  OAI22_X1 U2134 ( .A1(n18864), .A2(n18943), .B1(n1252), .B2(n18280), .ZN(
        n3706) );
  OAI22_X1 U2135 ( .A1(n18864), .A2(n18946), .B1(n1252), .B2(n18281), .ZN(
        n3707) );
  OAI22_X1 U2136 ( .A1(n18864), .A2(n18949), .B1(n18860), .B2(n18282), .ZN(
        n3708) );
  OAI22_X1 U2137 ( .A1(n18863), .A2(n18952), .B1(n18860), .B2(n18283), .ZN(
        n3709) );
  OAI22_X1 U2138 ( .A1(n18863), .A2(n18955), .B1(n18860), .B2(n18284), .ZN(
        n3710) );
  OAI22_X1 U2139 ( .A1(n18863), .A2(n18958), .B1(n18860), .B2(n18285), .ZN(
        n3711) );
  OAI22_X1 U2140 ( .A1(n1174), .A2(n18872), .B1(n18871), .B2(n17979), .ZN(
        n3720) );
  OAI22_X1 U2141 ( .A1(n1209), .A2(n18872), .B1(n18871), .B2(n17980), .ZN(
        n3721) );
  OAI22_X1 U2142 ( .A1(n18873), .A2(n18904), .B1(n18871), .B2(n17981), .ZN(
        n3725) );
  OAI22_X1 U2143 ( .A1(n18873), .A2(n18907), .B1(n18871), .B2(n17982), .ZN(
        n3726) );
  OAI22_X1 U2144 ( .A1(n18873), .A2(n18910), .B1(n18871), .B2(n17983), .ZN(
        n3727) );
  OAI22_X1 U2145 ( .A1(n18874), .A2(n18913), .B1(n18871), .B2(n17984), .ZN(
        n3728) );
  OAI22_X1 U2146 ( .A1(n18874), .A2(n18916), .B1(n18871), .B2(n17985), .ZN(
        n3729) );
  OAI22_X1 U2147 ( .A1(n18874), .A2(n18919), .B1(n18871), .B2(n17986), .ZN(
        n3730) );
  OAI22_X1 U2148 ( .A1(n18874), .A2(n18922), .B1(n18871), .B2(n17987), .ZN(
        n3731) );
  OAI22_X1 U2149 ( .A1(n18875), .A2(n18925), .B1(n1214), .B2(n17988), .ZN(
        n3732) );
  OAI22_X1 U2150 ( .A1(n18875), .A2(n18928), .B1(n1214), .B2(n17989), .ZN(
        n3733) );
  OAI22_X1 U2151 ( .A1(n18875), .A2(n18931), .B1(n1214), .B2(n17990), .ZN(
        n3734) );
  OAI22_X1 U2152 ( .A1(n18875), .A2(n18934), .B1(n1214), .B2(n17991), .ZN(
        n3735) );
  OAI22_X1 U2153 ( .A1(n18876), .A2(n18937), .B1(n1214), .B2(n17992), .ZN(
        n3736) );
  OAI22_X1 U2154 ( .A1(n18876), .A2(n18940), .B1(n1214), .B2(n17993), .ZN(
        n3737) );
  OAI22_X1 U2155 ( .A1(n18876), .A2(n18943), .B1(n1214), .B2(n17994), .ZN(
        n3738) );
  OAI22_X1 U2156 ( .A1(n18876), .A2(n18946), .B1(n18871), .B2(n17995), .ZN(
        n3739) );
  OAI22_X1 U2157 ( .A1(n18877), .A2(n18949), .B1(n18871), .B2(n17996), .ZN(
        n3740) );
  OAI22_X1 U2158 ( .A1(n18877), .A2(n18952), .B1(n18871), .B2(n17997), .ZN(
        n3741) );
  OAI22_X1 U2159 ( .A1(n18877), .A2(n18955), .B1(n18871), .B2(n17998), .ZN(
        n3742) );
  OAI22_X1 U2160 ( .A1(n18877), .A2(n18958), .B1(n18871), .B2(n17999), .ZN(
        n3743) );
  OAI22_X1 U2161 ( .A1(n1209), .A2(n18883), .B1(n18882), .B2(n17467), .ZN(
        n3753) );
  OAI22_X1 U2162 ( .A1(n18890), .A2(n18904), .B1(n18882), .B2(n17468), .ZN(
        n3757) );
  OAI22_X1 U2163 ( .A1(n18889), .A2(n18907), .B1(n18882), .B2(n17469), .ZN(
        n3758) );
  OAI22_X1 U2164 ( .A1(n18889), .A2(n18910), .B1(n18882), .B2(n17470), .ZN(
        n3759) );
  OAI22_X1 U2165 ( .A1(n18889), .A2(n18913), .B1(n18882), .B2(n17471), .ZN(
        n3760) );
  OAI22_X1 U2166 ( .A1(n18889), .A2(n18916), .B1(n18882), .B2(n17472), .ZN(
        n3761) );
  OAI22_X1 U2167 ( .A1(n18888), .A2(n18919), .B1(n18882), .B2(n17473), .ZN(
        n3762) );
  OAI22_X1 U2168 ( .A1(n18888), .A2(n18922), .B1(n18882), .B2(n17474), .ZN(
        n3763) );
  OAI22_X1 U2169 ( .A1(n18888), .A2(n18925), .B1(n1178), .B2(n17475), .ZN(
        n3764) );
  OAI22_X1 U2170 ( .A1(n18888), .A2(n18928), .B1(n1178), .B2(n17476), .ZN(
        n3765) );
  OAI22_X1 U2171 ( .A1(n18887), .A2(n18931), .B1(n1178), .B2(n17477), .ZN(
        n3766) );
  OAI22_X1 U2172 ( .A1(n18887), .A2(n18934), .B1(n1178), .B2(n17478), .ZN(
        n3767) );
  OAI22_X1 U2173 ( .A1(n18887), .A2(n18937), .B1(n1178), .B2(n17479), .ZN(
        n3768) );
  OAI22_X1 U2174 ( .A1(n18886), .A2(n18940), .B1(n1178), .B2(n17480), .ZN(
        n3769) );
  OAI22_X1 U2175 ( .A1(n18886), .A2(n18943), .B1(n1178), .B2(n17481), .ZN(
        n3770) );
  OAI22_X1 U2176 ( .A1(n18886), .A2(n18946), .B1(n18882), .B2(n17482), .ZN(
        n3771) );
  OAI22_X1 U2177 ( .A1(n18886), .A2(n18949), .B1(n18882), .B2(n17483), .ZN(
        n3772) );
  OAI22_X1 U2178 ( .A1(n18885), .A2(n18952), .B1(n18882), .B2(n17484), .ZN(
        n3773) );
  OAI22_X1 U2179 ( .A1(n18885), .A2(n18955), .B1(n18882), .B2(n17485), .ZN(
        n3774) );
  OAI22_X1 U2180 ( .A1(n18885), .A2(n18958), .B1(n18882), .B2(n17486), .ZN(
        n3775) );
  OAI22_X1 U2181 ( .A1(n1174), .A2(n18894), .B1(n18893), .B2(n17715), .ZN(
        n3784) );
  OAI22_X1 U2182 ( .A1(n18895), .A2(n18904), .B1(n18893), .B2(n17716), .ZN(
        n3789) );
  OAI22_X1 U2183 ( .A1(n18895), .A2(n18907), .B1(n18893), .B2(n17717), .ZN(
        n3790) );
  OAI22_X1 U2184 ( .A1(n18895), .A2(n18910), .B1(n18893), .B2(n17718), .ZN(
        n3791) );
  OAI22_X1 U2185 ( .A1(n18896), .A2(n18913), .B1(n18893), .B2(n17727), .ZN(
        n3792) );
  OAI22_X1 U2186 ( .A1(n18896), .A2(n18916), .B1(n18893), .B2(n17728), .ZN(
        n3793) );
  OAI22_X1 U2187 ( .A1(n18896), .A2(n18919), .B1(n18893), .B2(n17729), .ZN(
        n3794) );
  OAI22_X1 U2188 ( .A1(n18896), .A2(n18922), .B1(n18893), .B2(n17730), .ZN(
        n3795) );
  OAI22_X1 U2189 ( .A1(n18897), .A2(n18925), .B1(n1142), .B2(n17731), .ZN(
        n3796) );
  OAI22_X1 U2190 ( .A1(n18897), .A2(n18928), .B1(n1142), .B2(n17732), .ZN(
        n3797) );
  OAI22_X1 U2191 ( .A1(n18897), .A2(n18931), .B1(n1142), .B2(n17733), .ZN(
        n3798) );
  OAI22_X1 U2192 ( .A1(n18897), .A2(n18934), .B1(n1142), .B2(n17734), .ZN(
        n3799) );
  OAI22_X1 U2193 ( .A1(n18898), .A2(n18937), .B1(n1142), .B2(n17735), .ZN(
        n3800) );
  OAI22_X1 U2194 ( .A1(n18898), .A2(n18940), .B1(n1142), .B2(n17736), .ZN(
        n3801) );
  OAI22_X1 U2195 ( .A1(n18898), .A2(n18943), .B1(n1142), .B2(n17737), .ZN(
        n3802) );
  OAI22_X1 U2196 ( .A1(n18898), .A2(n18946), .B1(n18893), .B2(n17738), .ZN(
        n3803) );
  OAI22_X1 U2197 ( .A1(n18899), .A2(n18949), .B1(n18893), .B2(n17739), .ZN(
        n3804) );
  OAI22_X1 U2198 ( .A1(n18899), .A2(n18952), .B1(n18893), .B2(n17740), .ZN(
        n3805) );
  OAI22_X1 U2199 ( .A1(n18899), .A2(n18955), .B1(n18893), .B2(n17741), .ZN(
        n3806) );
  OAI22_X1 U2200 ( .A1(n18899), .A2(n18958), .B1(n18893), .B2(n17742), .ZN(
        n3807) );
  OAI21_X1 U2201 ( .B1(n1212), .B2(n2112), .A(n18999), .ZN(n2150) );
  OAI21_X1 U2202 ( .B1(n1176), .B2(n2112), .A(n18997), .ZN(n2116) );
  OAI21_X1 U2203 ( .B1(n1247), .B2(n1975), .A(n18999), .ZN(n2045) );
  OAI21_X1 U2204 ( .B1(n1247), .B2(n1838), .A(n18999), .ZN(n1908) );
  OAI21_X1 U2205 ( .B1(n1247), .B2(n1561), .A(n18998), .ZN(n1631) );
  OAI22_X1 U2206 ( .A1(n1209), .A2(n18561), .B1(n18570), .B2(n17495), .ZN(
        n2857) );
  OAI22_X1 U2207 ( .A1(n1282), .A2(n18561), .B1(n18570), .B2(n17496), .ZN(
        n2858) );
  OAI22_X1 U2208 ( .A1(n1419), .A2(n18561), .B1(n18570), .B2(n17497), .ZN(
        n2859) );
  OAI22_X1 U2209 ( .A1(n1694), .A2(n18561), .B1(n18569), .B2(n17498), .ZN(
        n2860) );
  OAI22_X1 U2210 ( .A1(n18561), .A2(n18906), .B1(n18569), .B2(n17499), .ZN(
        n2861) );
  OAI22_X1 U2211 ( .A1(n18562), .A2(n18909), .B1(n18569), .B2(n17500), .ZN(
        n2862) );
  OAI22_X1 U2212 ( .A1(n18561), .A2(n18912), .B1(n18569), .B2(n17501), .ZN(
        n2863) );
  OAI22_X1 U2213 ( .A1(n18562), .A2(n18915), .B1(n18568), .B2(n17502), .ZN(
        n2864) );
  OAI22_X1 U2214 ( .A1(n18561), .A2(n18918), .B1(n18568), .B2(n17503), .ZN(
        n2865) );
  OAI22_X1 U2215 ( .A1(n18562), .A2(n18921), .B1(n18568), .B2(n17504), .ZN(
        n2866) );
  OAI22_X1 U2216 ( .A1(n18561), .A2(n18924), .B1(n18568), .B2(n17505), .ZN(
        n2867) );
  OAI22_X1 U2217 ( .A1(n18562), .A2(n18927), .B1(n18567), .B2(n17506), .ZN(
        n2868) );
  OAI22_X1 U2218 ( .A1(n18562), .A2(n18930), .B1(n18567), .B2(n17507), .ZN(
        n2869) );
  OAI22_X1 U2219 ( .A1(n18562), .A2(n18933), .B1(n18567), .B2(n17508), .ZN(
        n2870) );
  OAI22_X1 U2220 ( .A1(n18562), .A2(n18936), .B1(n18567), .B2(n17509), .ZN(
        n2871) );
  OAI22_X1 U2221 ( .A1(n18562), .A2(n18939), .B1(n18566), .B2(n17510), .ZN(
        n2872) );
  OAI22_X1 U2222 ( .A1(n18562), .A2(n18942), .B1(n18566), .B2(n17511), .ZN(
        n2873) );
  OAI22_X1 U2223 ( .A1(n18562), .A2(n18945), .B1(n18566), .B2(n17512), .ZN(
        n2874) );
  OAI22_X1 U2224 ( .A1(n18562), .A2(n18948), .B1(n18566), .B2(n17513), .ZN(
        n2875) );
  OAI22_X1 U2225 ( .A1(n18562), .A2(n18951), .B1(n18565), .B2(n17514), .ZN(
        n2876) );
  OAI22_X1 U2226 ( .A1(n18562), .A2(n18954), .B1(n18565), .B2(n17515), .ZN(
        n2877) );
  OAI22_X1 U2227 ( .A1(n18562), .A2(n18957), .B1(n18565), .B2(n17516), .ZN(
        n2878) );
  OAI22_X1 U2228 ( .A1(n18562), .A2(n18960), .B1(n18565), .B2(n17517), .ZN(
        n2879) );
  OAI22_X1 U2229 ( .A1(n18561), .A2(n18963), .B1(n18564), .B2(n17487), .ZN(
        n2880) );
  OAI22_X1 U2230 ( .A1(n18561), .A2(n18966), .B1(n18564), .B2(n17488), .ZN(
        n2881) );
  OAI22_X1 U2231 ( .A1(n18561), .A2(n18969), .B1(n18564), .B2(n17489), .ZN(
        n2882) );
  OAI22_X1 U2232 ( .A1(n18561), .A2(n18972), .B1(n18564), .B2(n17490), .ZN(
        n2883) );
  OAI22_X1 U2233 ( .A1(n18561), .A2(n18975), .B1(n18563), .B2(n17491), .ZN(
        n2884) );
  OAI22_X1 U2234 ( .A1(n18561), .A2(n18978), .B1(n18563), .B2(n17492), .ZN(
        n2885) );
  OAI22_X1 U2235 ( .A1(n18561), .A2(n18981), .B1(n18563), .B2(n17493), .ZN(
        n2886) );
  OAI22_X1 U2236 ( .A1(n18562), .A2(n18993), .B1(n18563), .B2(n17494), .ZN(
        n2887) );
  OAI22_X1 U2237 ( .A1(n1174), .A2(n18575), .B1(n18584), .B2(n17583), .ZN(
        n2888) );
  OAI22_X1 U2238 ( .A1(n1282), .A2(n18575), .B1(n18584), .B2(n17584), .ZN(
        n2890) );
  OAI22_X1 U2239 ( .A1(n1419), .A2(n18575), .B1(n18584), .B2(n17585), .ZN(
        n2891) );
  OAI22_X1 U2240 ( .A1(n1694), .A2(n18575), .B1(n18583), .B2(n17586), .ZN(
        n2892) );
  OAI22_X1 U2241 ( .A1(n18575), .A2(n18906), .B1(n18583), .B2(n17587), .ZN(
        n2893) );
  OAI22_X1 U2242 ( .A1(n18576), .A2(n18909), .B1(n18583), .B2(n17588), .ZN(
        n2894) );
  OAI22_X1 U2243 ( .A1(n18575), .A2(n18912), .B1(n18583), .B2(n17589), .ZN(
        n2895) );
  OAI22_X1 U2244 ( .A1(n18576), .A2(n18915), .B1(n18582), .B2(n17590), .ZN(
        n2896) );
  OAI22_X1 U2245 ( .A1(n18575), .A2(n18918), .B1(n18582), .B2(n17591), .ZN(
        n2897) );
  OAI22_X1 U2246 ( .A1(n18576), .A2(n18921), .B1(n18582), .B2(n17592), .ZN(
        n2898) );
  OAI22_X1 U2247 ( .A1(n18575), .A2(n18924), .B1(n18582), .B2(n17593), .ZN(
        n2899) );
  OAI22_X1 U2248 ( .A1(n18576), .A2(n18927), .B1(n18581), .B2(n17594), .ZN(
        n2900) );
  OAI22_X1 U2249 ( .A1(n18576), .A2(n18930), .B1(n18581), .B2(n17595), .ZN(
        n2901) );
  OAI22_X1 U2250 ( .A1(n18576), .A2(n18933), .B1(n18581), .B2(n17596), .ZN(
        n2902) );
  OAI22_X1 U2251 ( .A1(n18576), .A2(n18936), .B1(n18580), .B2(n17597), .ZN(
        n2903) );
  OAI22_X1 U2252 ( .A1(n18576), .A2(n18939), .B1(n18580), .B2(n17598), .ZN(
        n2904) );
  OAI22_X1 U2253 ( .A1(n18576), .A2(n18942), .B1(n18580), .B2(n17599), .ZN(
        n2905) );
  OAI22_X1 U2254 ( .A1(n18576), .A2(n18945), .B1(n18580), .B2(n17600), .ZN(
        n2906) );
  OAI22_X1 U2255 ( .A1(n18576), .A2(n18948), .B1(n18579), .B2(n17601), .ZN(
        n2907) );
  OAI22_X1 U2256 ( .A1(n18576), .A2(n18951), .B1(n18579), .B2(n17602), .ZN(
        n2908) );
  OAI22_X1 U2257 ( .A1(n18576), .A2(n18954), .B1(n18579), .B2(n17603), .ZN(
        n2909) );
  OAI22_X1 U2258 ( .A1(n18576), .A2(n18957), .B1(n18579), .B2(n17604), .ZN(
        n2910) );
  OAI22_X1 U2259 ( .A1(n18576), .A2(n18960), .B1(n18578), .B2(n17605), .ZN(
        n2911) );
  OAI22_X1 U2260 ( .A1(n18575), .A2(n18963), .B1(n18578), .B2(n17606), .ZN(
        n2912) );
  OAI22_X1 U2261 ( .A1(n18575), .A2(n18966), .B1(n18578), .B2(n17607), .ZN(
        n2913) );
  OAI22_X1 U2262 ( .A1(n18575), .A2(n18969), .B1(n18578), .B2(n17608), .ZN(
        n2914) );
  OAI22_X1 U2263 ( .A1(n18575), .A2(n18972), .B1(n18577), .B2(n17609), .ZN(
        n2915) );
  OAI22_X1 U2264 ( .A1(n18575), .A2(n18975), .B1(n18577), .B2(n17610), .ZN(
        n2916) );
  OAI22_X1 U2265 ( .A1(n18575), .A2(n18978), .B1(n18577), .B2(n17611), .ZN(
        n2917) );
  OAI22_X1 U2266 ( .A1(n18575), .A2(n18981), .B1(n18577), .B2(n17612), .ZN(
        n2918) );
  OAI22_X1 U2267 ( .A1(n18576), .A2(n18993), .B1(n18581), .B2(n17613), .ZN(
        n2919) );
  OAI22_X1 U2268 ( .A1(n1174), .A2(n18601), .B1(n18610), .B2(n17638), .ZN(
        n2952) );
  OAI22_X1 U2269 ( .A1(n1209), .A2(n18601), .B1(n18610), .B2(n17639), .ZN(
        n2953) );
  OAI22_X1 U2270 ( .A1(n1419), .A2(n18601), .B1(n18610), .B2(n17640), .ZN(
        n2955) );
  OAI22_X1 U2271 ( .A1(n1694), .A2(n18601), .B1(n18609), .B2(n17641), .ZN(
        n2956) );
  OAI22_X1 U2272 ( .A1(n18601), .A2(n18906), .B1(n18609), .B2(n17642), .ZN(
        n2957) );
  OAI22_X1 U2273 ( .A1(n18602), .A2(n18909), .B1(n18609), .B2(n17643), .ZN(
        n2958) );
  OAI22_X1 U2274 ( .A1(n18601), .A2(n18912), .B1(n18609), .B2(n17644), .ZN(
        n2959) );
  OAI22_X1 U2275 ( .A1(n18602), .A2(n18915), .B1(n18608), .B2(n17645), .ZN(
        n2960) );
  OAI22_X1 U2276 ( .A1(n18601), .A2(n18918), .B1(n18608), .B2(n17646), .ZN(
        n2961) );
  OAI22_X1 U2277 ( .A1(n18602), .A2(n18921), .B1(n18608), .B2(n17647), .ZN(
        n2962) );
  OAI22_X1 U2278 ( .A1(n18601), .A2(n18924), .B1(n18608), .B2(n17648), .ZN(
        n2963) );
  OAI22_X1 U2279 ( .A1(n18602), .A2(n18927), .B1(n18607), .B2(n17649), .ZN(
        n2964) );
  OAI22_X1 U2280 ( .A1(n18602), .A2(n18930), .B1(n18607), .B2(n17650), .ZN(
        n2965) );
  OAI22_X1 U2281 ( .A1(n18602), .A2(n18933), .B1(n18607), .B2(n17651), .ZN(
        n2966) );
  OAI22_X1 U2282 ( .A1(n18602), .A2(n18936), .B1(n18606), .B2(n17652), .ZN(
        n2967) );
  OAI22_X1 U2283 ( .A1(n18602), .A2(n18939), .B1(n18606), .B2(n17653), .ZN(
        n2968) );
  OAI22_X1 U2284 ( .A1(n18602), .A2(n18942), .B1(n18606), .B2(n17654), .ZN(
        n2969) );
  OAI22_X1 U2285 ( .A1(n18602), .A2(n18945), .B1(n18606), .B2(n17655), .ZN(
        n2970) );
  OAI22_X1 U2286 ( .A1(n18602), .A2(n18948), .B1(n18605), .B2(n17656), .ZN(
        n2971) );
  OAI22_X1 U2287 ( .A1(n18602), .A2(n18951), .B1(n18605), .B2(n17657), .ZN(
        n2972) );
  OAI22_X1 U2288 ( .A1(n18602), .A2(n18954), .B1(n18605), .B2(n17658), .ZN(
        n2973) );
  OAI22_X1 U2289 ( .A1(n18602), .A2(n18957), .B1(n18605), .B2(n17659), .ZN(
        n2974) );
  OAI22_X1 U2290 ( .A1(n18602), .A2(n18960), .B1(n18604), .B2(n17660), .ZN(
        n2975) );
  OAI22_X1 U2291 ( .A1(n18601), .A2(n18963), .B1(n18604), .B2(n17661), .ZN(
        n2976) );
  OAI22_X1 U2292 ( .A1(n18601), .A2(n18966), .B1(n18604), .B2(n17662), .ZN(
        n2977) );
  OAI22_X1 U2293 ( .A1(n18601), .A2(n18969), .B1(n18604), .B2(n17663), .ZN(
        n2978) );
  OAI22_X1 U2294 ( .A1(n18601), .A2(n18972), .B1(n18603), .B2(n17664), .ZN(
        n2979) );
  OAI22_X1 U2295 ( .A1(n18601), .A2(n18975), .B1(n18603), .B2(n17665), .ZN(
        n2980) );
  OAI22_X1 U2296 ( .A1(n18601), .A2(n18978), .B1(n18603), .B2(n17666), .ZN(
        n2981) );
  OAI22_X1 U2297 ( .A1(n18601), .A2(n18981), .B1(n18603), .B2(n17667), .ZN(
        n2982) );
  OAI22_X1 U2298 ( .A1(n18602), .A2(n18993), .B1(n18607), .B2(n17668), .ZN(
        n2983) );
  OAI22_X1 U2299 ( .A1(n1174), .A2(n18648), .B1(n18657), .B2(n18192), .ZN(
        n3080) );
  OAI22_X1 U2300 ( .A1(n1209), .A2(n18648), .B1(n18657), .B2(n18193), .ZN(
        n3081) );
  OAI22_X1 U2301 ( .A1(n1282), .A2(n18648), .B1(n18657), .B2(n18194), .ZN(
        n3082) );
  OAI22_X1 U2302 ( .A1(n1694), .A2(n18648), .B1(n18656), .B2(n18195), .ZN(
        n3084) );
  OAI22_X1 U2303 ( .A1(n18648), .A2(n18905), .B1(n18656), .B2(n18196), .ZN(
        n3085) );
  OAI22_X1 U2304 ( .A1(n18649), .A2(n18908), .B1(n18656), .B2(n18197), .ZN(
        n3086) );
  OAI22_X1 U2305 ( .A1(n18648), .A2(n18911), .B1(n18656), .B2(n18198), .ZN(
        n3087) );
  OAI22_X1 U2306 ( .A1(n18649), .A2(n18914), .B1(n18655), .B2(n18199), .ZN(
        n3088) );
  OAI22_X1 U2307 ( .A1(n18648), .A2(n18917), .B1(n18655), .B2(n18200), .ZN(
        n3089) );
  OAI22_X1 U2308 ( .A1(n18649), .A2(n18920), .B1(n18655), .B2(n18201), .ZN(
        n3090) );
  OAI22_X1 U2309 ( .A1(n18648), .A2(n18923), .B1(n18655), .B2(n18202), .ZN(
        n3091) );
  OAI22_X1 U2310 ( .A1(n18649), .A2(n18926), .B1(n18654), .B2(n18203), .ZN(
        n3092) );
  OAI22_X1 U2311 ( .A1(n18649), .A2(n18929), .B1(n18654), .B2(n18204), .ZN(
        n3093) );
  OAI22_X1 U2312 ( .A1(n18649), .A2(n18932), .B1(n18654), .B2(n18205), .ZN(
        n3094) );
  OAI22_X1 U2313 ( .A1(n18649), .A2(n18935), .B1(n18653), .B2(n18206), .ZN(
        n3095) );
  OAI22_X1 U2314 ( .A1(n18649), .A2(n18938), .B1(n18653), .B2(n18207), .ZN(
        n3096) );
  OAI22_X1 U2315 ( .A1(n18649), .A2(n18941), .B1(n18653), .B2(n18208), .ZN(
        n3097) );
  OAI22_X1 U2316 ( .A1(n18649), .A2(n18944), .B1(n18653), .B2(n18209), .ZN(
        n3098) );
  OAI22_X1 U2317 ( .A1(n18649), .A2(n18947), .B1(n18652), .B2(n18210), .ZN(
        n3099) );
  OAI22_X1 U2318 ( .A1(n18649), .A2(n18950), .B1(n18652), .B2(n18211), .ZN(
        n3100) );
  OAI22_X1 U2319 ( .A1(n18649), .A2(n18953), .B1(n18652), .B2(n18212), .ZN(
        n3101) );
  OAI22_X1 U2320 ( .A1(n18649), .A2(n18956), .B1(n18652), .B2(n18213), .ZN(
        n3102) );
  OAI22_X1 U2321 ( .A1(n18649), .A2(n18959), .B1(n18651), .B2(n18214), .ZN(
        n3103) );
  OAI22_X1 U2322 ( .A1(n18648), .A2(n18962), .B1(n18651), .B2(n18215), .ZN(
        n3104) );
  OAI22_X1 U2323 ( .A1(n18648), .A2(n18965), .B1(n18651), .B2(n18216), .ZN(
        n3105) );
  OAI22_X1 U2324 ( .A1(n18648), .A2(n18968), .B1(n18651), .B2(n18217), .ZN(
        n3106) );
  OAI22_X1 U2325 ( .A1(n18648), .A2(n18971), .B1(n18650), .B2(n18218), .ZN(
        n3107) );
  OAI22_X1 U2326 ( .A1(n18648), .A2(n18974), .B1(n18650), .B2(n18219), .ZN(
        n3108) );
  OAI22_X1 U2327 ( .A1(n18648), .A2(n18977), .B1(n18650), .B2(n18220), .ZN(
        n3109) );
  OAI22_X1 U2328 ( .A1(n18648), .A2(n18980), .B1(n18650), .B2(n18221), .ZN(
        n3110) );
  OAI22_X1 U2329 ( .A1(n18649), .A2(n18992), .B1(n18654), .B2(n18222), .ZN(
        n3111) );
  OAI22_X1 U2330 ( .A1(n1174), .A2(n18739), .B1(n18748), .B2(n18223), .ZN(
        n3336) );
  OAI22_X1 U2331 ( .A1(n1209), .A2(n18739), .B1(n18748), .B2(n18224), .ZN(
        n3337) );
  OAI22_X1 U2332 ( .A1(n1282), .A2(n18739), .B1(n18748), .B2(n18225), .ZN(
        n3338) );
  OAI22_X1 U2333 ( .A1(n1419), .A2(n18739), .B1(n18747), .B2(n18226), .ZN(
        n3339) );
  OAI22_X1 U2334 ( .A1(n18739), .A2(n18905), .B1(n18747), .B2(n18227), .ZN(
        n3341) );
  OAI22_X1 U2335 ( .A1(n18739), .A2(n18908), .B1(n18747), .B2(n18228), .ZN(
        n3342) );
  OAI22_X1 U2336 ( .A1(n18739), .A2(n18911), .B1(n18747), .B2(n18229), .ZN(
        n3343) );
  OAI22_X1 U2337 ( .A1(n18739), .A2(n18914), .B1(n18746), .B2(n18238), .ZN(
        n3344) );
  OAI22_X1 U2338 ( .A1(n18739), .A2(n18917), .B1(n18746), .B2(n18239), .ZN(
        n3345) );
  OAI22_X1 U2339 ( .A1(n18739), .A2(n18920), .B1(n18746), .B2(n18240), .ZN(
        n3346) );
  OAI22_X1 U2340 ( .A1(n18739), .A2(n18923), .B1(n18746), .B2(n18241), .ZN(
        n3347) );
  OAI22_X1 U2341 ( .A1(n18739), .A2(n18926), .B1(n18745), .B2(n18242), .ZN(
        n3348) );
  OAI22_X1 U2342 ( .A1(n18740), .A2(n18929), .B1(n18745), .B2(n18243), .ZN(
        n3349) );
  OAI22_X1 U2343 ( .A1(n18740), .A2(n18932), .B1(n18745), .B2(n18244), .ZN(
        n3350) );
  OAI22_X1 U2344 ( .A1(n18740), .A2(n18935), .B1(n18744), .B2(n18245), .ZN(
        n3351) );
  OAI22_X1 U2345 ( .A1(n18740), .A2(n18938), .B1(n18744), .B2(n18246), .ZN(
        n3352) );
  OAI22_X1 U2346 ( .A1(n18740), .A2(n18941), .B1(n18744), .B2(n18247), .ZN(
        n3353) );
  OAI22_X1 U2347 ( .A1(n18740), .A2(n18944), .B1(n18744), .B2(n18248), .ZN(
        n3354) );
  OAI22_X1 U2348 ( .A1(n18740), .A2(n18947), .B1(n18743), .B2(n18249), .ZN(
        n3355) );
  OAI22_X1 U2349 ( .A1(n18740), .A2(n18950), .B1(n18743), .B2(n18250), .ZN(
        n3356) );
  OAI22_X1 U2350 ( .A1(n18740), .A2(n18953), .B1(n18743), .B2(n18251), .ZN(
        n3357) );
  OAI22_X1 U2351 ( .A1(n18740), .A2(n18956), .B1(n18743), .B2(n18252), .ZN(
        n3358) );
  OAI22_X1 U2352 ( .A1(n18740), .A2(n18959), .B1(n18742), .B2(n18253), .ZN(
        n3359) );
  OAI22_X1 U2353 ( .A1(n18740), .A2(n18962), .B1(n18742), .B2(n18230), .ZN(
        n3360) );
  OAI22_X1 U2354 ( .A1(n18740), .A2(n18965), .B1(n18742), .B2(n18231), .ZN(
        n3361) );
  OAI22_X1 U2355 ( .A1(n18740), .A2(n18968), .B1(n18742), .B2(n18232), .ZN(
        n3362) );
  OAI22_X1 U2356 ( .A1(n18739), .A2(n18971), .B1(n18741), .B2(n18233), .ZN(
        n3363) );
  OAI22_X1 U2357 ( .A1(n18740), .A2(n18974), .B1(n18741), .B2(n18234), .ZN(
        n3364) );
  OAI22_X1 U2358 ( .A1(n18739), .A2(n18977), .B1(n18741), .B2(n18235), .ZN(
        n3365) );
  OAI22_X1 U2359 ( .A1(n18740), .A2(n18980), .B1(n18741), .B2(n18236), .ZN(
        n3366) );
  OAI22_X1 U2360 ( .A1(n18739), .A2(n18992), .B1(n18745), .B2(n18237), .ZN(
        n3367) );
  BUF_X1 U2361 ( .A(RESET), .Z(n18996) );
  OAI21_X1 U2362 ( .B1(n1138), .B2(n1247), .A(n18997), .ZN(n1214) );
  OAI21_X1 U2363 ( .B1(n1138), .B2(n1212), .A(n18997), .ZN(n1178) );
  OAI21_X1 U2364 ( .B1(n1138), .B2(n1176), .A(n18997), .ZN(n1142) );
  OAI21_X1 U2365 ( .B1(n1139), .B2(n2112), .A(n18997), .ZN(n2079) );
  OAI21_X1 U2366 ( .B1(n1212), .B2(n1975), .A(n18999), .ZN(n2011) );
  OAI21_X1 U2367 ( .B1(n1176), .B2(n1975), .A(n18999), .ZN(n1977) );
  OAI21_X1 U2368 ( .B1(n1139), .B2(n1975), .A(n18999), .ZN(n1942) );
  OAI21_X1 U2369 ( .B1(n1212), .B2(n1838), .A(n18999), .ZN(n1874) );
  OAI21_X1 U2370 ( .B1(n1176), .B2(n1838), .A(n18999), .ZN(n1840) );
  OAI21_X1 U2371 ( .B1(n1139), .B2(n1838), .A(n18999), .ZN(n1805) );
  OAI21_X1 U2372 ( .B1(n1247), .B2(n1700), .A(n18999), .ZN(n1770) );
  OAI21_X1 U2373 ( .B1(n1212), .B2(n1700), .A(n18999), .ZN(n1736) );
  OAI21_X1 U2374 ( .B1(n1176), .B2(n1700), .A(n18999), .ZN(n1702) );
  OAI21_X1 U2375 ( .B1(n1212), .B2(n1561), .A(n18998), .ZN(n1597) );
  OAI21_X1 U2376 ( .B1(n1176), .B2(n1561), .A(n18998), .ZN(n1563) );
  OAI21_X1 U2377 ( .B1(n1139), .B2(n1561), .A(n18998), .ZN(n1528) );
  OAI21_X1 U2378 ( .B1(n1247), .B2(n1424), .A(n18998), .ZN(n1494) );
  OAI21_X1 U2379 ( .B1(n1212), .B2(n1424), .A(n18998), .ZN(n1460) );
  OAI21_X1 U2380 ( .B1(n1176), .B2(n1424), .A(n18998), .ZN(n1426) );
  OAI21_X1 U2381 ( .B1(n1139), .B2(n1424), .A(n18998), .ZN(n1390) );
  OAI21_X1 U2382 ( .B1(n1247), .B2(n1286), .A(n18998), .ZN(n1356) );
  OAI21_X1 U2383 ( .B1(n1212), .B2(n1286), .A(n18998), .ZN(n1322) );
  OAI21_X1 U2384 ( .B1(n1176), .B2(n1286), .A(n18998), .ZN(n1288) );
  OAI21_X1 U2385 ( .B1(n1139), .B2(n1286), .A(n18998), .ZN(n1252) );
  NAND2_X1 U2386 ( .A1(n2113), .A2(n2114), .ZN(n1139) );
  OAI221_X1 U2387 ( .B1(n17383), .B2(n18546), .C1(n17669), .C2(n18543), .A(
        n3904), .ZN(n3903) );
  AOI22_X1 U2388 ( .A1(n18540), .A2(net535500), .B1(n18538), .B2(OUT1[0]), 
        .ZN(n3904) );
  OAI221_X1 U2389 ( .B1(n17384), .B2(n18546), .C1(n17670), .C2(n18543), .A(
        n3885), .ZN(n3884) );
  AOI22_X1 U2390 ( .A1(n18540), .A2(net535501), .B1(n18538), .B2(OUT1[1]), 
        .ZN(n3885) );
  OAI221_X1 U2391 ( .B1(n17385), .B2(n18546), .C1(n17671), .C2(n18543), .A(
        n3866), .ZN(n3865) );
  AOI22_X1 U2392 ( .A1(n18540), .A2(net535502), .B1(n18539), .B2(OUT1[2]), 
        .ZN(n3866) );
  OAI221_X1 U2393 ( .B1(n17386), .B2(n18546), .C1(n17672), .C2(n18543), .A(
        n2759), .ZN(n2758) );
  AOI22_X1 U2394 ( .A1(n18540), .A2(net535503), .B1(n18538), .B2(OUT1[3]), 
        .ZN(n2759) );
  OAI221_X1 U2395 ( .B1(n17387), .B2(n18546), .C1(n17673), .C2(n18543), .A(
        n2740), .ZN(n2739) );
  AOI22_X1 U2396 ( .A1(n18540), .A2(net535504), .B1(n18538), .B2(OUT1[4]), 
        .ZN(n2740) );
  OAI221_X1 U2397 ( .B1(n17388), .B2(n18546), .C1(n17674), .C2(n18543), .A(
        n2721), .ZN(n2720) );
  AOI22_X1 U2398 ( .A1(n18540), .A2(net535505), .B1(n18538), .B2(OUT1[5]), 
        .ZN(n2721) );
  OAI221_X1 U2399 ( .B1(n17389), .B2(n18546), .C1(n17675), .C2(n18543), .A(
        n2702), .ZN(n2701) );
  AOI22_X1 U2400 ( .A1(n18540), .A2(net535506), .B1(n18538), .B2(OUT1[6]), 
        .ZN(n2702) );
  OAI221_X1 U2401 ( .B1(n17390), .B2(n18546), .C1(n17676), .C2(n18543), .A(
        n2683), .ZN(n2682) );
  AOI22_X1 U2402 ( .A1(n18540), .A2(net535507), .B1(n18538), .B2(OUT1[7]), 
        .ZN(n2683) );
  OAI221_X1 U2403 ( .B1(n17719), .B2(n18537), .C1(n18230), .C2(n18534), .A(
        n2361), .ZN(n2358) );
  AOI22_X1 U2404 ( .A1(n18531), .A2(net366975), .B1(n18526), .B2(net310782), 
        .ZN(n2361) );
  OAI221_X1 U2405 ( .B1(n17720), .B2(n18537), .C1(n18231), .C2(n18534), .A(
        n2342), .ZN(n2339) );
  AOI22_X1 U2406 ( .A1(n18531), .A2(net366976), .B1(n18526), .B2(net310783), 
        .ZN(n2342) );
  OAI221_X1 U2407 ( .B1(n17721), .B2(n18537), .C1(n18232), .C2(n18534), .A(
        n2323), .ZN(n2320) );
  AOI22_X1 U2408 ( .A1(n18531), .A2(net366977), .B1(n18526), .B2(net310784), 
        .ZN(n2323) );
  OAI221_X1 U2409 ( .B1(n17722), .B2(n18537), .C1(n18233), .C2(n18534), .A(
        n2304), .ZN(n2301) );
  AOI22_X1 U2410 ( .A1(n18531), .A2(net366978), .B1(n18526), .B2(net310785), 
        .ZN(n2304) );
  OAI221_X1 U2411 ( .B1(n17723), .B2(n18537), .C1(n18234), .C2(n18534), .A(
        n2285), .ZN(n2282) );
  AOI22_X1 U2412 ( .A1(n18531), .A2(net366979), .B1(n18526), .B2(net310786), 
        .ZN(n2285) );
  OAI221_X1 U2413 ( .B1(n17724), .B2(n18537), .C1(n18235), .C2(n18534), .A(
        n2266), .ZN(n2263) );
  AOI22_X1 U2414 ( .A1(n18531), .A2(net366980), .B1(n18526), .B2(net310787), 
        .ZN(n2266) );
  OAI221_X1 U2415 ( .B1(n17725), .B2(n18537), .C1(n18236), .C2(n18534), .A(
        n2247), .ZN(n2244) );
  AOI22_X1 U2416 ( .A1(n18531), .A2(net366981), .B1(n18526), .B2(net310788), 
        .ZN(n2247) );
  OAI221_X1 U2417 ( .B1(n17726), .B2(n18537), .C1(n18237), .C2(n18534), .A(
        n2201), .ZN(n2192) );
  AOI22_X1 U2418 ( .A1(n18531), .A2(net366982), .B1(n18526), .B2(net310789), 
        .ZN(n2201) );
  OAI221_X1 U2419 ( .B1(n17727), .B2(n18535), .C1(n18238), .C2(n18532), .A(
        n2665), .ZN(n2662) );
  AOI22_X1 U2420 ( .A1(n18529), .A2(net366959), .B1(n18527), .B2(net310766), 
        .ZN(n2665) );
  OAI221_X1 U2421 ( .B1(n17728), .B2(n18535), .C1(n18239), .C2(n18532), .A(
        n2646), .ZN(n2643) );
  AOI22_X1 U2422 ( .A1(n18529), .A2(net366960), .B1(n18527), .B2(net310767), 
        .ZN(n2646) );
  OAI221_X1 U2423 ( .B1(n17729), .B2(n18535), .C1(n18240), .C2(n18532), .A(
        n2627), .ZN(n2624) );
  AOI22_X1 U2424 ( .A1(n18529), .A2(net366961), .B1(n18527), .B2(net310768), 
        .ZN(n2627) );
  OAI221_X1 U2425 ( .B1(n17730), .B2(n18535), .C1(n18241), .C2(n18532), .A(
        n2608), .ZN(n2605) );
  AOI22_X1 U2426 ( .A1(n18529), .A2(net366962), .B1(n18527), .B2(net310769), 
        .ZN(n2608) );
  OAI221_X1 U2427 ( .B1(n17731), .B2(n18536), .C1(n18242), .C2(n18533), .A(
        n2589), .ZN(n2586) );
  AOI22_X1 U2428 ( .A1(n18530), .A2(net366963), .B1(n18527), .B2(net310770), 
        .ZN(n2589) );
  OAI221_X1 U2429 ( .B1(n17732), .B2(n18536), .C1(n18243), .C2(n18533), .A(
        n2570), .ZN(n2567) );
  AOI22_X1 U2430 ( .A1(n18530), .A2(net366964), .B1(n18527), .B2(net310771), 
        .ZN(n2570) );
  OAI221_X1 U2431 ( .B1(n17733), .B2(n18536), .C1(n18244), .C2(n18533), .A(
        n2551), .ZN(n2548) );
  AOI22_X1 U2432 ( .A1(n18530), .A2(net366965), .B1(n18527), .B2(net310772), 
        .ZN(n2551) );
  OAI221_X1 U2433 ( .B1(n17734), .B2(n18536), .C1(n18245), .C2(n18533), .A(
        n2532), .ZN(n2529) );
  AOI22_X1 U2434 ( .A1(n18530), .A2(net366966), .B1(n18527), .B2(net310773), 
        .ZN(n2532) );
  OAI221_X1 U2435 ( .B1(n17735), .B2(n18536), .C1(n18246), .C2(n18533), .A(
        n2513), .ZN(n2510) );
  AOI22_X1 U2436 ( .A1(n18530), .A2(net366967), .B1(n18527), .B2(net310774), 
        .ZN(n2513) );
  OAI221_X1 U2437 ( .B1(n17736), .B2(n18536), .C1(n18247), .C2(n18533), .A(
        n2494), .ZN(n2491) );
  AOI22_X1 U2438 ( .A1(n18530), .A2(net366968), .B1(n18527), .B2(net310775), 
        .ZN(n2494) );
  OAI221_X1 U2439 ( .B1(n17737), .B2(n18536), .C1(n18248), .C2(n18533), .A(
        n2475), .ZN(n2472) );
  AOI22_X1 U2440 ( .A1(n18530), .A2(net366969), .B1(n18527), .B2(net310776), 
        .ZN(n2475) );
  OAI221_X1 U2441 ( .B1(n17738), .B2(n18536), .C1(n18249), .C2(n18533), .A(
        n2456), .ZN(n2453) );
  AOI22_X1 U2442 ( .A1(n18530), .A2(net366970), .B1(n18527), .B2(net310777), 
        .ZN(n2456) );
  OAI221_X1 U2443 ( .B1(n17739), .B2(n18536), .C1(n18250), .C2(n18533), .A(
        n2437), .ZN(n2434) );
  AOI22_X1 U2444 ( .A1(n18530), .A2(net366971), .B1(n18526), .B2(net310778), 
        .ZN(n2437) );
  OAI221_X1 U2445 ( .B1(n17740), .B2(n18536), .C1(n18251), .C2(n18533), .A(
        n2418), .ZN(n2415) );
  AOI22_X1 U2446 ( .A1(n18530), .A2(net366972), .B1(n18526), .B2(net310779), 
        .ZN(n2418) );
  OAI221_X1 U2447 ( .B1(n17741), .B2(n18536), .C1(n18252), .C2(n18533), .A(
        n2399), .ZN(n2396) );
  AOI22_X1 U2448 ( .A1(n18530), .A2(net366973), .B1(n18526), .B2(net310780), 
        .ZN(n2399) );
  OAI221_X1 U2449 ( .B1(n17742), .B2(n18536), .C1(n18253), .C2(n18533), .A(
        n2380), .ZN(n2377) );
  AOI22_X1 U2450 ( .A1(n18530), .A2(net366974), .B1(n18526), .B2(net310781), 
        .ZN(n2380) );
  OAI221_X1 U2451 ( .B1(n17487), .B2(n18415), .C1(n17840), .C2(n18412), .A(
        n4101), .ZN(n4094) );
  AOI22_X1 U2452 ( .A1(n18409), .A2(net423198), .B1(n18404), .B2(net591747), 
        .ZN(n4101) );
  OAI221_X1 U2453 ( .B1(n17488), .B2(n18415), .C1(n17841), .C2(n18412), .A(
        n4083), .ZN(n4076) );
  AOI22_X1 U2454 ( .A1(n18409), .A2(net423199), .B1(n18404), .B2(net591748), 
        .ZN(n4083) );
  OAI221_X1 U2455 ( .B1(n17489), .B2(n18415), .C1(n17842), .C2(n18412), .A(
        n4065), .ZN(n4058) );
  AOI22_X1 U2456 ( .A1(n18409), .A2(net423200), .B1(n18404), .B2(net591749), 
        .ZN(n4065) );
  OAI221_X1 U2457 ( .B1(n17490), .B2(n18415), .C1(n17843), .C2(n18412), .A(
        n4047), .ZN(n4040) );
  AOI22_X1 U2458 ( .A1(n18409), .A2(net423201), .B1(n18404), .B2(net591750), 
        .ZN(n4047) );
  OAI221_X1 U2459 ( .B1(n17491), .B2(n18415), .C1(n17844), .C2(n18412), .A(
        n4029), .ZN(n4022) );
  AOI22_X1 U2460 ( .A1(n18409), .A2(net423202), .B1(n18404), .B2(net591751), 
        .ZN(n4029) );
  OAI221_X1 U2461 ( .B1(n17492), .B2(n18415), .C1(n17845), .C2(n18412), .A(
        n4011), .ZN(n4004) );
  AOI22_X1 U2462 ( .A1(n18409), .A2(net423203), .B1(n18404), .B2(net591752), 
        .ZN(n4011) );
  OAI221_X1 U2463 ( .B1(n17493), .B2(n18415), .C1(n17846), .C2(n18412), .A(
        n3993), .ZN(n3986) );
  AOI22_X1 U2464 ( .A1(n18409), .A2(net423204), .B1(n18404), .B2(net591753), 
        .ZN(n3993) );
  OAI221_X1 U2465 ( .B1(n17494), .B2(n18415), .C1(n17847), .C2(n18412), .A(
        n3956), .ZN(n3935) );
  AOI22_X1 U2466 ( .A1(n18409), .A2(net423205), .B1(n18404), .B2(net591754), 
        .ZN(n3956) );
  OAI221_X1 U2467 ( .B1(n17518), .B2(n18413), .C1(n17848), .C2(n18410), .A(
        n4544), .ZN(n4526) );
  AOI22_X1 U2468 ( .A1(n18407), .A2(net423174), .B1(n18406), .B2(net591723), 
        .ZN(n4544) );
  OAI221_X1 U2469 ( .B1(n17495), .B2(n18413), .C1(n17849), .C2(n18410), .A(
        n4515), .ZN(n4508) );
  AOI22_X1 U2470 ( .A1(n18407), .A2(net423175), .B1(n18406), .B2(net591724), 
        .ZN(n4515) );
  OAI221_X1 U2471 ( .B1(n17496), .B2(n18413), .C1(n17850), .C2(n18410), .A(
        n4497), .ZN(n4490) );
  AOI22_X1 U2472 ( .A1(n18407), .A2(net423176), .B1(n18406), .B2(net591725), 
        .ZN(n4497) );
  OAI221_X1 U2473 ( .B1(n17497), .B2(n18413), .C1(n17851), .C2(n18410), .A(
        n4479), .ZN(n4472) );
  AOI22_X1 U2474 ( .A1(n18407), .A2(net423177), .B1(n18406), .B2(net591726), 
        .ZN(n4479) );
  OAI221_X1 U2475 ( .B1(n17498), .B2(n18413), .C1(n17852), .C2(n18410), .A(
        n4461), .ZN(n4454) );
  AOI22_X1 U2476 ( .A1(n18407), .A2(net423178), .B1(n18406), .B2(net591727), 
        .ZN(n4461) );
  OAI221_X1 U2477 ( .B1(n17499), .B2(n18413), .C1(n17853), .C2(n18410), .A(
        n4443), .ZN(n4436) );
  AOI22_X1 U2478 ( .A1(n18407), .A2(net423179), .B1(n18406), .B2(net591728), 
        .ZN(n4443) );
  OAI221_X1 U2479 ( .B1(n17500), .B2(n18413), .C1(n17854), .C2(n18410), .A(
        n4425), .ZN(n4418) );
  AOI22_X1 U2480 ( .A1(n18407), .A2(net423180), .B1(n18406), .B2(net591729), 
        .ZN(n4425) );
  OAI221_X1 U2481 ( .B1(n17501), .B2(n18413), .C1(n17855), .C2(n18410), .A(
        n4407), .ZN(n4400) );
  AOI22_X1 U2482 ( .A1(n18407), .A2(net423181), .B1(n18406), .B2(net591730), 
        .ZN(n4407) );
  OAI221_X1 U2483 ( .B1(n17502), .B2(n18413), .C1(n17856), .C2(n18410), .A(
        n4389), .ZN(n4382) );
  AOI22_X1 U2484 ( .A1(n18407), .A2(net423182), .B1(n18405), .B2(net591731), 
        .ZN(n4389) );
  OAI221_X1 U2485 ( .B1(n17503), .B2(n18413), .C1(n17857), .C2(n18410), .A(
        n4371), .ZN(n4364) );
  AOI22_X1 U2486 ( .A1(n18407), .A2(net423183), .B1(n18405), .B2(net591732), 
        .ZN(n4371) );
  OAI221_X1 U2487 ( .B1(n17504), .B2(n18413), .C1(n17858), .C2(n18410), .A(
        n4353), .ZN(n4346) );
  AOI22_X1 U2488 ( .A1(n18407), .A2(net423184), .B1(n18405), .B2(net591733), 
        .ZN(n4353) );
  OAI221_X1 U2489 ( .B1(n17505), .B2(n18413), .C1(n17859), .C2(n18410), .A(
        n4335), .ZN(n4328) );
  AOI22_X1 U2490 ( .A1(n18407), .A2(net423185), .B1(n18405), .B2(net591734), 
        .ZN(n4335) );
  OAI221_X1 U2491 ( .B1(n17506), .B2(n18414), .C1(n17860), .C2(n18411), .A(
        n4317), .ZN(n4310) );
  AOI22_X1 U2492 ( .A1(n18408), .A2(net423186), .B1(n18405), .B2(net591735), 
        .ZN(n4317) );
  OAI221_X1 U2493 ( .B1(n17507), .B2(n18414), .C1(n17861), .C2(n18411), .A(
        n4299), .ZN(n4292) );
  AOI22_X1 U2494 ( .A1(n18408), .A2(net423187), .B1(n18405), .B2(net591736), 
        .ZN(n4299) );
  OAI221_X1 U2495 ( .B1(n17508), .B2(n18414), .C1(n17862), .C2(n18411), .A(
        n4281), .ZN(n4274) );
  AOI22_X1 U2496 ( .A1(n18408), .A2(net423188), .B1(n18405), .B2(net591737), 
        .ZN(n4281) );
  OAI221_X1 U2497 ( .B1(n17509), .B2(n18414), .C1(n17863), .C2(n18411), .A(
        n4263), .ZN(n4256) );
  AOI22_X1 U2498 ( .A1(n18408), .A2(net423189), .B1(n18405), .B2(net591738), 
        .ZN(n4263) );
  OAI221_X1 U2499 ( .B1(n17510), .B2(n18414), .C1(n17864), .C2(n18411), .A(
        n4245), .ZN(n4238) );
  AOI22_X1 U2500 ( .A1(n18408), .A2(net423190), .B1(n18405), .B2(net591739), 
        .ZN(n4245) );
  OAI221_X1 U2501 ( .B1(n17511), .B2(n18414), .C1(n17865), .C2(n18411), .A(
        n4227), .ZN(n4220) );
  AOI22_X1 U2502 ( .A1(n18408), .A2(net423191), .B1(n18405), .B2(net591740), 
        .ZN(n4227) );
  OAI221_X1 U2503 ( .B1(n17512), .B2(n18414), .C1(n17866), .C2(n18411), .A(
        n4209), .ZN(n4202) );
  AOI22_X1 U2504 ( .A1(n18408), .A2(net423192), .B1(n18405), .B2(net591741), 
        .ZN(n4209) );
  OAI221_X1 U2505 ( .B1(n17513), .B2(n18414), .C1(n17867), .C2(n18411), .A(
        n4191), .ZN(n4184) );
  AOI22_X1 U2506 ( .A1(n18408), .A2(net423193), .B1(n18405), .B2(net591742), 
        .ZN(n4191) );
  OAI221_X1 U2507 ( .B1(n17514), .B2(n18414), .C1(n17868), .C2(n18411), .A(
        n4173), .ZN(n4166) );
  AOI22_X1 U2508 ( .A1(n18408), .A2(net423194), .B1(n18404), .B2(net591743), 
        .ZN(n4173) );
  OAI221_X1 U2509 ( .B1(n17515), .B2(n18414), .C1(n17869), .C2(n18411), .A(
        n4155), .ZN(n4148) );
  AOI22_X1 U2510 ( .A1(n18408), .A2(net423195), .B1(n18404), .B2(net591744), 
        .ZN(n4155) );
  OAI221_X1 U2511 ( .B1(n17516), .B2(n18414), .C1(n17870), .C2(n18411), .A(
        n4137), .ZN(n4130) );
  AOI22_X1 U2512 ( .A1(n18408), .A2(net423196), .B1(n18404), .B2(net591745), 
        .ZN(n4137) );
  OAI221_X1 U2513 ( .B1(n17517), .B2(n18414), .C1(n17871), .C2(n18411), .A(
        n4119), .ZN(n4112) );
  AOI22_X1 U2514 ( .A1(n18408), .A2(net423197), .B1(n18404), .B2(net591746), 
        .ZN(n4119) );
  AOI22_X1 U2515 ( .A1(n18507), .A2(net479401), .B1(net591555), .B2(n18504), 
        .ZN(n2363) );
  AOI22_X1 U2516 ( .A1(n18507), .A2(net479402), .B1(net591556), .B2(n18504), 
        .ZN(n2344) );
  AOI22_X1 U2517 ( .A1(n18507), .A2(net479403), .B1(net591557), .B2(n18504), 
        .ZN(n2325) );
  AOI22_X1 U2518 ( .A1(n18507), .A2(net479404), .B1(net591558), .B2(n18504), 
        .ZN(n2306) );
  AOI22_X1 U2519 ( .A1(n18507), .A2(net479405), .B1(net591559), .B2(n18504), 
        .ZN(n2287) );
  AOI22_X1 U2520 ( .A1(n18507), .A2(net479406), .B1(net591560), .B2(n18504), 
        .ZN(n2268) );
  AOI22_X1 U2521 ( .A1(n18507), .A2(net479407), .B1(net591561), .B2(n18504), 
        .ZN(n2249) );
  AOI22_X1 U2522 ( .A1(n18442), .A2(net367111), .B1(n18440), .B2(OUT2[0]), 
        .ZN(n4530) );
  AOI22_X1 U2523 ( .A1(n18442), .A2(net367112), .B1(n18441), .B2(OUT2[1]), 
        .ZN(n4512) );
  AOI22_X1 U2524 ( .A1(n18442), .A2(net367113), .B1(n18441), .B2(OUT2[2]), 
        .ZN(n4494) );
  AOI22_X1 U2525 ( .A1(n18442), .A2(net367114), .B1(n18441), .B2(OUT2[3]), 
        .ZN(n4476) );
  AOI22_X1 U2526 ( .A1(n18442), .A2(net367115), .B1(n18441), .B2(OUT2[4]), 
        .ZN(n4458) );
  AOI22_X1 U2527 ( .A1(n18442), .A2(net367116), .B1(n18441), .B2(OUT2[5]), 
        .ZN(n4440) );
  AOI22_X1 U2528 ( .A1(n18442), .A2(net367117), .B1(n18441), .B2(OUT2[6]), 
        .ZN(n4422) );
  AOI22_X1 U2529 ( .A1(n18442), .A2(net367118), .B1(n18441), .B2(OUT2[7]), 
        .ZN(n4404) );
  AOI22_X1 U2530 ( .A1(n18442), .A2(net367119), .B1(n18441), .B2(OUT2[8]), 
        .ZN(n4386) );
  AOI22_X1 U2531 ( .A1(n18442), .A2(net367120), .B1(n18440), .B2(OUT2[9]), 
        .ZN(n4368) );
  AOI22_X1 U2532 ( .A1(n18442), .A2(net367121), .B1(n18440), .B2(OUT2[10]), 
        .ZN(n4350) );
  AOI22_X1 U2533 ( .A1(n18442), .A2(net367122), .B1(n18440), .B2(OUT2[11]), 
        .ZN(n4332) );
  AOI22_X1 U2534 ( .A1(n18443), .A2(net367123), .B1(n18440), .B2(OUT2[12]), 
        .ZN(n4314) );
  AOI22_X1 U2535 ( .A1(n18443), .A2(net367124), .B1(n18440), .B2(OUT2[13]), 
        .ZN(n4296) );
  AOI22_X1 U2536 ( .A1(n18443), .A2(net367125), .B1(n18440), .B2(OUT2[14]), 
        .ZN(n4278) );
  AOI22_X1 U2537 ( .A1(n18443), .A2(net367126), .B1(n18440), .B2(OUT2[15]), 
        .ZN(n4260) );
  AOI22_X1 U2538 ( .A1(n18443), .A2(net367127), .B1(n18440), .B2(OUT2[16]), 
        .ZN(n4242) );
  AOI22_X1 U2539 ( .A1(n18443), .A2(net367128), .B1(n18440), .B2(OUT2[17]), 
        .ZN(n4224) );
  AOI22_X1 U2540 ( .A1(n18443), .A2(net367129), .B1(n18440), .B2(OUT2[18]), 
        .ZN(n4206) );
  AOI22_X1 U2541 ( .A1(n18443), .A2(net367130), .B1(n18440), .B2(OUT2[19]), 
        .ZN(n4188) );
  AOI22_X1 U2542 ( .A1(n18443), .A2(net367131), .B1(n18440), .B2(OUT2[20]), 
        .ZN(n4170) );
  AOI22_X1 U2543 ( .A1(n18443), .A2(net367132), .B1(n18440), .B2(OUT2[21]), 
        .ZN(n4152) );
  AOI22_X1 U2544 ( .A1(n18443), .A2(net367133), .B1(n18440), .B2(OUT2[22]), 
        .ZN(n4134) );
  AOI22_X1 U2545 ( .A1(n18443), .A2(net367134), .B1(n18440), .B2(OUT2[23]), 
        .ZN(n4116) );
  AOI22_X1 U2546 ( .A1(n18444), .A2(net367135), .B1(n18440), .B2(OUT2[24]), 
        .ZN(n4098) );
  AOI22_X1 U2547 ( .A1(n18444), .A2(net367136), .B1(n18440), .B2(OUT2[25]), 
        .ZN(n4080) );
  AOI22_X1 U2548 ( .A1(n18444), .A2(net367137), .B1(n18440), .B2(OUT2[26]), 
        .ZN(n4062) );
  AOI22_X1 U2549 ( .A1(n18444), .A2(net367138), .B1(n18440), .B2(OUT2[27]), 
        .ZN(n4044) );
  AOI22_X1 U2550 ( .A1(n18444), .A2(net367139), .B1(n18440), .B2(OUT2[28]), 
        .ZN(n4026) );
  AOI22_X1 U2551 ( .A1(n18444), .A2(net367140), .B1(n18440), .B2(OUT2[29]), 
        .ZN(n4008) );
  AOI22_X1 U2552 ( .A1(n18444), .A2(net367141), .B1(n18440), .B2(OUT2[30]), 
        .ZN(n3990) );
  AOI22_X1 U2553 ( .A1(n18444), .A2(net367142), .B1(n18440), .B2(OUT2[31]), 
        .ZN(n3941) );
  AOI22_X1 U2554 ( .A1(n18529), .A2(net366951), .B1(n18528), .B2(net310758), 
        .ZN(n3910) );
  AOI22_X1 U2555 ( .A1(n18517), .A2(net591659), .B1(n18516), .B2(net591627), 
        .ZN(n3916) );
  AOI22_X1 U2556 ( .A1(n18529), .A2(net366952), .B1(n18528), .B2(net310759), 
        .ZN(n3886) );
  AOI22_X1 U2557 ( .A1(n18517), .A2(net591660), .B1(n18516), .B2(net591628), 
        .ZN(n3887) );
  AOI22_X1 U2558 ( .A1(n18529), .A2(net366953), .B1(n18528), .B2(net310760), 
        .ZN(n3867) );
  AOI22_X1 U2559 ( .A1(n18517), .A2(net591661), .B1(n18516), .B2(net591629), 
        .ZN(n3868) );
  AOI22_X1 U2560 ( .A1(n18529), .A2(net366954), .B1(n18528), .B2(net310761), 
        .ZN(n3848) );
  AOI22_X1 U2561 ( .A1(n18517), .A2(net591662), .B1(n18516), .B2(net591630), 
        .ZN(n3849) );
  AOI22_X1 U2562 ( .A1(n18529), .A2(net366955), .B1(n18528), .B2(net310762), 
        .ZN(n2741) );
  AOI22_X1 U2563 ( .A1(n18517), .A2(net591663), .B1(n18516), .B2(net591631), 
        .ZN(n2742) );
  AOI22_X1 U2564 ( .A1(n18529), .A2(net366956), .B1(n18528), .B2(net310763), 
        .ZN(n2722) );
  AOI22_X1 U2565 ( .A1(n18517), .A2(net591664), .B1(n18516), .B2(net591632), 
        .ZN(n2723) );
  AOI22_X1 U2566 ( .A1(n18529), .A2(net366957), .B1(n18528), .B2(net310764), 
        .ZN(n2703) );
  AOI22_X1 U2567 ( .A1(n18517), .A2(net591665), .B1(n18516), .B2(net591633), 
        .ZN(n2704) );
  AOI22_X1 U2568 ( .A1(n18529), .A2(net366958), .B1(n18528), .B2(net310765), 
        .ZN(n2684) );
  AOI22_X1 U2569 ( .A1(n18517), .A2(net591666), .B1(n18516), .B2(net591634), 
        .ZN(n2685) );
  AOI22_X1 U2570 ( .A1(n18540), .A2(net535508), .B1(n18538), .B2(OUT1[8]), 
        .ZN(n2664) );
  AOI22_X1 U2571 ( .A1(n18517), .A2(net591667), .B1(n18515), .B2(net591635), 
        .ZN(n2666) );
  AOI22_X1 U2572 ( .A1(n18540), .A2(net535509), .B1(n18539), .B2(OUT1[9]), 
        .ZN(n2645) );
  AOI22_X1 U2573 ( .A1(n18517), .A2(net591668), .B1(n18515), .B2(net591636), 
        .ZN(n2647) );
  AOI22_X1 U2574 ( .A1(n18540), .A2(net535510), .B1(n18538), .B2(OUT1[10]), 
        .ZN(n2626) );
  AOI22_X1 U2575 ( .A1(n18517), .A2(net591669), .B1(n18515), .B2(net591637), 
        .ZN(n2628) );
  AOI22_X1 U2576 ( .A1(n18540), .A2(net535511), .B1(n18538), .B2(OUT1[11]), 
        .ZN(n2607) );
  AOI22_X1 U2577 ( .A1(n18517), .A2(net591670), .B1(n18515), .B2(net591638), 
        .ZN(n2609) );
  AOI22_X1 U2578 ( .A1(n18541), .A2(net535512), .B1(n18538), .B2(OUT1[12]), 
        .ZN(n2588) );
  AOI22_X1 U2579 ( .A1(n18518), .A2(net591671), .B1(n18515), .B2(net591639), 
        .ZN(n2590) );
  AOI22_X1 U2580 ( .A1(n18541), .A2(net535513), .B1(n18538), .B2(OUT1[13]), 
        .ZN(n2569) );
  AOI22_X1 U2581 ( .A1(n18518), .A2(net591672), .B1(n18515), .B2(net591640), 
        .ZN(n2571) );
  AOI22_X1 U2582 ( .A1(n18541), .A2(net535514), .B1(n18538), .B2(OUT1[14]), 
        .ZN(n2550) );
  AOI22_X1 U2583 ( .A1(n18518), .A2(net591673), .B1(n18515), .B2(net591641), 
        .ZN(n2552) );
  AOI22_X1 U2584 ( .A1(n18541), .A2(net535515), .B1(n18538), .B2(OUT1[15]), 
        .ZN(n2531) );
  AOI22_X1 U2585 ( .A1(n18518), .A2(net591674), .B1(n18515), .B2(net591642), 
        .ZN(n2533) );
  AOI22_X1 U2586 ( .A1(n18541), .A2(net535516), .B1(n18538), .B2(OUT1[16]), 
        .ZN(n2512) );
  AOI22_X1 U2587 ( .A1(n18518), .A2(net591675), .B1(n18515), .B2(net591643), 
        .ZN(n2514) );
  AOI22_X1 U2588 ( .A1(n18541), .A2(net535517), .B1(n18538), .B2(OUT1[17]), 
        .ZN(n2493) );
  AOI22_X1 U2589 ( .A1(n18518), .A2(net591676), .B1(n18515), .B2(net591644), 
        .ZN(n2495) );
  AOI22_X1 U2590 ( .A1(n18541), .A2(net535518), .B1(n18538), .B2(OUT1[18]), 
        .ZN(n2474) );
  AOI22_X1 U2591 ( .A1(n18518), .A2(net591677), .B1(n18515), .B2(net591645), 
        .ZN(n2476) );
  AOI22_X1 U2592 ( .A1(n18541), .A2(net535519), .B1(n18538), .B2(OUT1[19]), 
        .ZN(n2455) );
  AOI22_X1 U2593 ( .A1(n18518), .A2(net591678), .B1(n18515), .B2(net591646), 
        .ZN(n2457) );
  AOI22_X1 U2594 ( .A1(n18541), .A2(net535520), .B1(n18538), .B2(OUT1[20]), 
        .ZN(n2436) );
  AOI22_X1 U2595 ( .A1(n18518), .A2(net591679), .B1(n18514), .B2(net591647), 
        .ZN(n2438) );
  AOI22_X1 U2596 ( .A1(n18541), .A2(net535521), .B1(n18538), .B2(OUT1[21]), 
        .ZN(n2417) );
  AOI22_X1 U2597 ( .A1(n18518), .A2(net591680), .B1(n18514), .B2(net591648), 
        .ZN(n2419) );
  AOI22_X1 U2598 ( .A1(n18541), .A2(net535522), .B1(n18538), .B2(OUT1[22]), 
        .ZN(n2398) );
  AOI22_X1 U2599 ( .A1(n18518), .A2(net591681), .B1(n18514), .B2(net591649), 
        .ZN(n2400) );
  AOI22_X1 U2600 ( .A1(n18541), .A2(net535523), .B1(n18538), .B2(OUT1[23]), 
        .ZN(n2379) );
  AOI22_X1 U2601 ( .A1(n18518), .A2(net591682), .B1(n18514), .B2(net591650), 
        .ZN(n2381) );
  AOI22_X1 U2602 ( .A1(n18519), .A2(net591683), .B1(n18514), .B2(net591651), 
        .ZN(n2362) );
  AOI22_X1 U2603 ( .A1(n18542), .A2(net535524), .B1(n18539), .B2(OUT1[24]), 
        .ZN(n2360) );
  AOI22_X1 U2604 ( .A1(n18519), .A2(net591684), .B1(n18514), .B2(net591652), 
        .ZN(n2343) );
  AOI22_X1 U2605 ( .A1(n18542), .A2(net535525), .B1(n18539), .B2(OUT1[25]), 
        .ZN(n2341) );
  AOI22_X1 U2606 ( .A1(n18519), .A2(net591685), .B1(n18514), .B2(net591653), 
        .ZN(n2324) );
  AOI22_X1 U2607 ( .A1(n18542), .A2(net535526), .B1(n18539), .B2(OUT1[26]), 
        .ZN(n2322) );
  AOI22_X1 U2608 ( .A1(n18519), .A2(net591686), .B1(n18514), .B2(net591654), 
        .ZN(n2305) );
  AOI22_X1 U2609 ( .A1(n18542), .A2(net535527), .B1(n18539), .B2(OUT1[27]), 
        .ZN(n2303) );
  AOI22_X1 U2610 ( .A1(n18519), .A2(net591687), .B1(n18514), .B2(net591655), 
        .ZN(n2286) );
  AOI22_X1 U2611 ( .A1(n18542), .A2(net535528), .B1(n18539), .B2(OUT1[28]), 
        .ZN(n2284) );
  AOI22_X1 U2612 ( .A1(n18519), .A2(net591688), .B1(n18514), .B2(net591656), 
        .ZN(n2267) );
  AOI22_X1 U2613 ( .A1(n18542), .A2(net535529), .B1(n18539), .B2(OUT1[29]), 
        .ZN(n2265) );
  AOI22_X1 U2614 ( .A1(n18519), .A2(net591689), .B1(n18514), .B2(net591657), 
        .ZN(n2248) );
  AOI22_X1 U2615 ( .A1(n18542), .A2(net535530), .B1(n18539), .B2(OUT1[30]), 
        .ZN(n2246) );
  AOI22_X1 U2616 ( .A1(n18519), .A2(net591690), .B1(n18514), .B2(net591658), 
        .ZN(n2206) );
  AOI22_X1 U2617 ( .A1(n18542), .A2(net535531), .B1(n18539), .B2(OUT1[31]), 
        .ZN(n2196) );
  AOI22_X1 U2618 ( .A1(n18419), .A2(net367015), .B1(n18418), .B2(net479410), 
        .ZN(n4541) );
  AOI22_X1 U2619 ( .A1(n18431), .A2(net310502), .B1(n18430), .B2(net535436), 
        .ZN(n4536) );
  AOI22_X1 U2620 ( .A1(n18419), .A2(net367016), .B1(n18418), .B2(net479411), 
        .ZN(n4514) );
  AOI22_X1 U2621 ( .A1(n18431), .A2(net310503), .B1(n18430), .B2(net535437), 
        .ZN(n4513) );
  AOI22_X1 U2622 ( .A1(n18419), .A2(net367017), .B1(n18418), .B2(net479412), 
        .ZN(n4496) );
  AOI22_X1 U2623 ( .A1(n18431), .A2(net310504), .B1(n18430), .B2(net535438), 
        .ZN(n4495) );
  AOI22_X1 U2624 ( .A1(n18419), .A2(net367018), .B1(n18418), .B2(net479413), 
        .ZN(n4478) );
  AOI22_X1 U2625 ( .A1(n18431), .A2(net310505), .B1(n18430), .B2(net535439), 
        .ZN(n4477) );
  AOI22_X1 U2626 ( .A1(n18419), .A2(net367019), .B1(n18418), .B2(net479414), 
        .ZN(n4460) );
  AOI22_X1 U2627 ( .A1(n18431), .A2(net310506), .B1(n18430), .B2(net535440), 
        .ZN(n4459) );
  AOI22_X1 U2628 ( .A1(n18419), .A2(net367020), .B1(n18418), .B2(net479415), 
        .ZN(n4442) );
  AOI22_X1 U2629 ( .A1(n18431), .A2(net310507), .B1(n18430), .B2(net535441), 
        .ZN(n4441) );
  AOI22_X1 U2630 ( .A1(n18419), .A2(net367021), .B1(n18418), .B2(net479416), 
        .ZN(n4424) );
  AOI22_X1 U2631 ( .A1(n18431), .A2(net310508), .B1(n18430), .B2(net535442), 
        .ZN(n4423) );
  AOI22_X1 U2632 ( .A1(n18419), .A2(net367022), .B1(n18418), .B2(net479417), 
        .ZN(n4406) );
  AOI22_X1 U2633 ( .A1(n18431), .A2(net310509), .B1(n18430), .B2(net535443), 
        .ZN(n4405) );
  AOI22_X1 U2634 ( .A1(n18419), .A2(net367023), .B1(n18417), .B2(net479418), 
        .ZN(n4388) );
  AOI22_X1 U2635 ( .A1(n18431), .A2(net310510), .B1(n18429), .B2(net535444), 
        .ZN(n4387) );
  AOI22_X1 U2636 ( .A1(n18419), .A2(net367024), .B1(n18417), .B2(net479419), 
        .ZN(n4370) );
  AOI22_X1 U2637 ( .A1(n18431), .A2(net310511), .B1(n18429), .B2(net535445), 
        .ZN(n4369) );
  AOI22_X1 U2638 ( .A1(n18419), .A2(net367025), .B1(n18417), .B2(net479420), 
        .ZN(n4352) );
  AOI22_X1 U2639 ( .A1(n18431), .A2(net310512), .B1(n18429), .B2(net535446), 
        .ZN(n4351) );
  AOI22_X1 U2640 ( .A1(n18419), .A2(net367026), .B1(n18417), .B2(net479421), 
        .ZN(n4334) );
  AOI22_X1 U2641 ( .A1(n18431), .A2(net310513), .B1(n18429), .B2(net535447), 
        .ZN(n4333) );
  AOI22_X1 U2642 ( .A1(n18420), .A2(net367027), .B1(n18417), .B2(net479422), 
        .ZN(n4316) );
  AOI22_X1 U2643 ( .A1(n18432), .A2(net310514), .B1(n18429), .B2(net535448), 
        .ZN(n4315) );
  AOI22_X1 U2644 ( .A1(n18420), .A2(net367028), .B1(n18417), .B2(net479423), 
        .ZN(n4298) );
  AOI22_X1 U2645 ( .A1(n18432), .A2(net310515), .B1(n18429), .B2(net535449), 
        .ZN(n4297) );
  AOI22_X1 U2646 ( .A1(n18420), .A2(net367029), .B1(n18417), .B2(net479424), 
        .ZN(n4280) );
  AOI22_X1 U2647 ( .A1(n18432), .A2(net310516), .B1(n18429), .B2(net535450), 
        .ZN(n4279) );
  AOI22_X1 U2648 ( .A1(n18420), .A2(net367030), .B1(n18417), .B2(net479425), 
        .ZN(n4262) );
  AOI22_X1 U2649 ( .A1(n18432), .A2(net310517), .B1(n18429), .B2(net535451), 
        .ZN(n4261) );
  AOI22_X1 U2650 ( .A1(n18420), .A2(net367031), .B1(n18417), .B2(net479426), 
        .ZN(n4244) );
  AOI22_X1 U2651 ( .A1(n18432), .A2(net310518), .B1(n18429), .B2(net535452), 
        .ZN(n4243) );
  AOI22_X1 U2652 ( .A1(n18420), .A2(net367032), .B1(n18417), .B2(net479427), 
        .ZN(n4226) );
  AOI22_X1 U2653 ( .A1(n18432), .A2(net310519), .B1(n18429), .B2(net535453), 
        .ZN(n4225) );
  AOI22_X1 U2654 ( .A1(n18420), .A2(net367033), .B1(n18417), .B2(net479428), 
        .ZN(n4208) );
  AOI22_X1 U2655 ( .A1(n18432), .A2(net310520), .B1(n18429), .B2(net535454), 
        .ZN(n4207) );
  AOI22_X1 U2656 ( .A1(n18420), .A2(net367034), .B1(n18417), .B2(net479429), 
        .ZN(n4190) );
  AOI22_X1 U2657 ( .A1(n18432), .A2(net310521), .B1(n18429), .B2(net535455), 
        .ZN(n4189) );
  AOI22_X1 U2658 ( .A1(n18420), .A2(net367035), .B1(n18416), .B2(net479430), 
        .ZN(n4172) );
  AOI22_X1 U2659 ( .A1(n18432), .A2(net310522), .B1(n18428), .B2(net535456), 
        .ZN(n4171) );
  AOI22_X1 U2660 ( .A1(n18420), .A2(net367036), .B1(n18416), .B2(net479431), 
        .ZN(n4154) );
  AOI22_X1 U2661 ( .A1(n18432), .A2(net310523), .B1(n18428), .B2(net535457), 
        .ZN(n4153) );
  AOI22_X1 U2662 ( .A1(n18420), .A2(net367037), .B1(n18416), .B2(net479432), 
        .ZN(n4136) );
  AOI22_X1 U2663 ( .A1(n18432), .A2(net310524), .B1(n18428), .B2(net535458), 
        .ZN(n4135) );
  AOI22_X1 U2664 ( .A1(n18420), .A2(net367038), .B1(n18416), .B2(net479433), 
        .ZN(n4118) );
  AOI22_X1 U2665 ( .A1(n18432), .A2(net310525), .B1(n18428), .B2(net535459), 
        .ZN(n4117) );
  AOI22_X1 U2666 ( .A1(n18421), .A2(net367039), .B1(n18416), .B2(net479434), 
        .ZN(n4100) );
  AOI22_X1 U2667 ( .A1(n18433), .A2(net310526), .B1(n18428), .B2(net535460), 
        .ZN(n4099) );
  AOI22_X1 U2668 ( .A1(n18421), .A2(net367040), .B1(n18416), .B2(net479435), 
        .ZN(n4082) );
  AOI22_X1 U2669 ( .A1(n18433), .A2(net310527), .B1(n18428), .B2(net535461), 
        .ZN(n4081) );
  AOI22_X1 U2670 ( .A1(n18421), .A2(net367041), .B1(n18416), .B2(net479436), 
        .ZN(n4064) );
  AOI22_X1 U2671 ( .A1(n18433), .A2(net310528), .B1(n18428), .B2(net535462), 
        .ZN(n4063) );
  AOI22_X1 U2672 ( .A1(n18421), .A2(net367042), .B1(n18416), .B2(net479437), 
        .ZN(n4046) );
  AOI22_X1 U2673 ( .A1(n18433), .A2(net310529), .B1(n18428), .B2(net535463), 
        .ZN(n4045) );
  AOI22_X1 U2674 ( .A1(n18421), .A2(net367043), .B1(n18416), .B2(net479438), 
        .ZN(n4028) );
  AOI22_X1 U2675 ( .A1(n18433), .A2(net310530), .B1(n18428), .B2(net535464), 
        .ZN(n4027) );
  AOI22_X1 U2676 ( .A1(n18421), .A2(net367044), .B1(n18416), .B2(net479439), 
        .ZN(n4010) );
  AOI22_X1 U2677 ( .A1(n18433), .A2(net310531), .B1(n18428), .B2(net535465), 
        .ZN(n4009) );
  AOI22_X1 U2678 ( .A1(n18421), .A2(net367045), .B1(n18416), .B2(net479440), 
        .ZN(n3992) );
  AOI22_X1 U2679 ( .A1(n18433), .A2(net310532), .B1(n18428), .B2(net535466), 
        .ZN(n3991) );
  AOI22_X1 U2680 ( .A1(n18421), .A2(net367046), .B1(n18416), .B2(net479441), 
        .ZN(n3951) );
  AOI22_X1 U2681 ( .A1(n18433), .A2(net310533), .B1(n18428), .B2(net535467), 
        .ZN(n3946) );
  AOI22_X1 U2682 ( .A1(n18505), .A2(net479377), .B1(net591531), .B2(n18502), 
        .ZN(n3918) );
  AOI22_X1 U2683 ( .A1(n18505), .A2(net479378), .B1(net591532), .B2(n18502), 
        .ZN(n3888) );
  AOI22_X1 U2684 ( .A1(n18505), .A2(net479379), .B1(net591533), .B2(n18502), 
        .ZN(n3869) );
  AOI22_X1 U2685 ( .A1(n18505), .A2(net479380), .B1(net591534), .B2(n18502), 
        .ZN(n3850) );
  AOI22_X1 U2686 ( .A1(n18505), .A2(net479381), .B1(net591535), .B2(n18502), 
        .ZN(n2743) );
  AOI22_X1 U2687 ( .A1(n18505), .A2(net479382), .B1(net591536), .B2(n18502), 
        .ZN(n2724) );
  AOI22_X1 U2688 ( .A1(n18505), .A2(net479383), .B1(net591537), .B2(n18502), 
        .ZN(n2705) );
  AOI22_X1 U2689 ( .A1(n18505), .A2(net479384), .B1(net591538), .B2(n18502), 
        .ZN(n2686) );
  AOI22_X1 U2690 ( .A1(n18505), .A2(net479385), .B1(net591539), .B2(n18502), 
        .ZN(n2667) );
  AOI22_X1 U2691 ( .A1(n18505), .A2(net479386), .B1(net591540), .B2(n18502), 
        .ZN(n2648) );
  AOI22_X1 U2692 ( .A1(n18505), .A2(net479387), .B1(net591541), .B2(n18502), 
        .ZN(n2629) );
  AOI22_X1 U2693 ( .A1(n18505), .A2(net479388), .B1(net591542), .B2(n18502), 
        .ZN(n2610) );
  AOI22_X1 U2694 ( .A1(n18506), .A2(net479389), .B1(net591543), .B2(n18503), 
        .ZN(n2591) );
  AOI22_X1 U2695 ( .A1(n18506), .A2(net479390), .B1(net591544), .B2(n18503), 
        .ZN(n2572) );
  AOI22_X1 U2696 ( .A1(n18506), .A2(net479391), .B1(net591545), .B2(n18503), 
        .ZN(n2553) );
  AOI22_X1 U2697 ( .A1(n18506), .A2(net479392), .B1(net591546), .B2(n18503), 
        .ZN(n2534) );
  AOI22_X1 U2698 ( .A1(n18506), .A2(net479393), .B1(net591547), .B2(n18503), 
        .ZN(n2515) );
  AOI22_X1 U2699 ( .A1(n18506), .A2(net479394), .B1(net591548), .B2(n18503), 
        .ZN(n2496) );
  AOI22_X1 U2700 ( .A1(n18506), .A2(net479395), .B1(net591549), .B2(n18503), 
        .ZN(n2477) );
  AOI22_X1 U2701 ( .A1(n18506), .A2(net479396), .B1(net591550), .B2(n18503), 
        .ZN(n2458) );
  AOI22_X1 U2702 ( .A1(n18506), .A2(net479397), .B1(net591551), .B2(n18503), 
        .ZN(n2439) );
  AOI22_X1 U2703 ( .A1(n18506), .A2(net479398), .B1(net591552), .B2(n18503), 
        .ZN(n2420) );
  AOI22_X1 U2704 ( .A1(n18506), .A2(net479399), .B1(net591553), .B2(n18503), 
        .ZN(n2401) );
  AOI22_X1 U2705 ( .A1(n18506), .A2(net479400), .B1(net591554), .B2(n18503), 
        .ZN(n2382) );
  AOI22_X1 U2706 ( .A1(n18507), .A2(net479408), .B1(n18504), .B2(net591562), 
        .ZN(n2211) );
  NAND4_X1 U2707 ( .A1(n4522), .A2(n4523), .A3(n4524), .A4(n4525), .ZN(n2760)
         );
  AOI221_X1 U2708 ( .B1(n18362), .B2(net366951), .C1(n18359), .C2(net591787), 
        .A(n4555), .ZN(n4522) );
  NOR4_X1 U2709 ( .A1(n4546), .A2(n4547), .A3(n4548), .A4(n4549), .ZN(n4524)
         );
  AOI221_X1 U2710 ( .B1(n18374), .B2(net535468), .C1(n18371), .C2(net591531), 
        .A(n4554), .ZN(n4523) );
  NAND4_X1 U2711 ( .A1(n4504), .A2(n4505), .A3(n4506), .A4(n4507), .ZN(n2761)
         );
  AOI221_X1 U2712 ( .B1(n18362), .B2(net366952), .C1(n18359), .C2(net591788), 
        .A(n4521), .ZN(n4504) );
  NOR4_X1 U2713 ( .A1(n4516), .A2(n4517), .A3(n4518), .A4(n4519), .ZN(n4506)
         );
  AOI221_X1 U2714 ( .B1(n18374), .B2(net535469), .C1(n18371), .C2(net591532), 
        .A(n4520), .ZN(n4505) );
  NAND4_X1 U2715 ( .A1(n4486), .A2(n4487), .A3(n4488), .A4(n4489), .ZN(n2762)
         );
  AOI221_X1 U2716 ( .B1(n18362), .B2(net366953), .C1(n18359), .C2(net591789), 
        .A(n4503), .ZN(n4486) );
  NOR4_X1 U2717 ( .A1(n4498), .A2(n4499), .A3(n4500), .A4(n4501), .ZN(n4488)
         );
  AOI221_X1 U2718 ( .B1(n18374), .B2(net535470), .C1(n18371), .C2(net591533), 
        .A(n4502), .ZN(n4487) );
  NAND4_X1 U2719 ( .A1(n4468), .A2(n4469), .A3(n4470), .A4(n4471), .ZN(n2763)
         );
  AOI221_X1 U2720 ( .B1(n18362), .B2(net366954), .C1(n18359), .C2(net591790), 
        .A(n4485), .ZN(n4468) );
  NOR4_X1 U2721 ( .A1(n4480), .A2(n4481), .A3(n4482), .A4(n4483), .ZN(n4470)
         );
  AOI221_X1 U2722 ( .B1(n18374), .B2(net535471), .C1(n18371), .C2(net591534), 
        .A(n4484), .ZN(n4469) );
  NAND4_X1 U2723 ( .A1(n4450), .A2(n4451), .A3(n4452), .A4(n4453), .ZN(n2764)
         );
  AOI221_X1 U2724 ( .B1(n18362), .B2(net366955), .C1(n18359), .C2(net591791), 
        .A(n4467), .ZN(n4450) );
  NOR4_X1 U2725 ( .A1(n4462), .A2(n4463), .A3(n4464), .A4(n4465), .ZN(n4452)
         );
  AOI221_X1 U2726 ( .B1(n18374), .B2(net535472), .C1(n18371), .C2(net591535), 
        .A(n4466), .ZN(n4451) );
  NAND4_X1 U2727 ( .A1(n4432), .A2(n4433), .A3(n4434), .A4(n4435), .ZN(n2765)
         );
  AOI221_X1 U2728 ( .B1(n18362), .B2(net366956), .C1(n18359), .C2(net591792), 
        .A(n4449), .ZN(n4432) );
  NOR4_X1 U2729 ( .A1(n4444), .A2(n4445), .A3(n4446), .A4(n4447), .ZN(n4434)
         );
  AOI221_X1 U2730 ( .B1(n18374), .B2(net535473), .C1(n18371), .C2(net591536), 
        .A(n4448), .ZN(n4433) );
  NAND4_X1 U2731 ( .A1(n4414), .A2(n4415), .A3(n4416), .A4(n4417), .ZN(n2766)
         );
  AOI221_X1 U2732 ( .B1(n18362), .B2(net366957), .C1(n18359), .C2(net591793), 
        .A(n4431), .ZN(n4414) );
  NOR4_X1 U2733 ( .A1(n4426), .A2(n4427), .A3(n4428), .A4(n4429), .ZN(n4416)
         );
  AOI221_X1 U2734 ( .B1(n18374), .B2(net535474), .C1(n18371), .C2(net591537), 
        .A(n4430), .ZN(n4415) );
  NAND4_X1 U2735 ( .A1(n4396), .A2(n4397), .A3(n4398), .A4(n4399), .ZN(n2767)
         );
  AOI221_X1 U2736 ( .B1(n18362), .B2(net366958), .C1(n18359), .C2(net591794), 
        .A(n4413), .ZN(n4396) );
  NOR4_X1 U2737 ( .A1(n4408), .A2(n4409), .A3(n4410), .A4(n4411), .ZN(n4398)
         );
  AOI221_X1 U2738 ( .B1(n18374), .B2(net535475), .C1(n18371), .C2(net591538), 
        .A(n4412), .ZN(n4397) );
  NAND4_X1 U2739 ( .A1(n4378), .A2(n4379), .A3(n4380), .A4(n4381), .ZN(n2768)
         );
  AOI221_X1 U2740 ( .B1(n18362), .B2(net366959), .C1(n18359), .C2(net591795), 
        .A(n4395), .ZN(n4378) );
  NOR4_X1 U2741 ( .A1(n4390), .A2(n4391), .A3(n4392), .A4(n4393), .ZN(n4380)
         );
  AOI221_X1 U2742 ( .B1(n18374), .B2(net535476), .C1(n18371), .C2(net591539), 
        .A(n4394), .ZN(n4379) );
  NAND4_X1 U2743 ( .A1(n4360), .A2(n4361), .A3(n4362), .A4(n4363), .ZN(n2769)
         );
  AOI221_X1 U2744 ( .B1(n18362), .B2(net366960), .C1(n18359), .C2(net591796), 
        .A(n4377), .ZN(n4360) );
  NOR4_X1 U2745 ( .A1(n4372), .A2(n4373), .A3(n4374), .A4(n4375), .ZN(n4362)
         );
  AOI221_X1 U2746 ( .B1(n18374), .B2(net535477), .C1(n18371), .C2(net591540), 
        .A(n4376), .ZN(n4361) );
  NAND4_X1 U2747 ( .A1(n4342), .A2(n4343), .A3(n4344), .A4(n4345), .ZN(n2770)
         );
  AOI221_X1 U2748 ( .B1(n18362), .B2(net366961), .C1(n18359), .C2(net591797), 
        .A(n4359), .ZN(n4342) );
  NOR4_X1 U2749 ( .A1(n4354), .A2(n4355), .A3(n4356), .A4(n4357), .ZN(n4344)
         );
  AOI221_X1 U2750 ( .B1(n18374), .B2(net535478), .C1(n18371), .C2(net591541), 
        .A(n4358), .ZN(n4343) );
  NAND4_X1 U2751 ( .A1(n4324), .A2(n4325), .A3(n4326), .A4(n4327), .ZN(n2771)
         );
  AOI221_X1 U2752 ( .B1(n18362), .B2(net366962), .C1(n18359), .C2(net591798), 
        .A(n4341), .ZN(n4324) );
  NOR4_X1 U2753 ( .A1(n4336), .A2(n4337), .A3(n4338), .A4(n4339), .ZN(n4326)
         );
  AOI221_X1 U2754 ( .B1(n18374), .B2(net535479), .C1(n18371), .C2(net591542), 
        .A(n4340), .ZN(n4325) );
  NAND4_X1 U2755 ( .A1(n4306), .A2(n4307), .A3(n4308), .A4(n4309), .ZN(n2772)
         );
  AOI221_X1 U2756 ( .B1(n18363), .B2(net366963), .C1(n18360), .C2(net591799), 
        .A(n4323), .ZN(n4306) );
  NOR4_X1 U2757 ( .A1(n4318), .A2(n4319), .A3(n4320), .A4(n4321), .ZN(n4308)
         );
  AOI221_X1 U2758 ( .B1(n18375), .B2(net535480), .C1(n18372), .C2(net591543), 
        .A(n4322), .ZN(n4307) );
  NAND4_X1 U2759 ( .A1(n4288), .A2(n4289), .A3(n4290), .A4(n4291), .ZN(n2773)
         );
  AOI221_X1 U2760 ( .B1(n18363), .B2(net366964), .C1(n18360), .C2(net591800), 
        .A(n4305), .ZN(n4288) );
  NOR4_X1 U2761 ( .A1(n4300), .A2(n4301), .A3(n4302), .A4(n4303), .ZN(n4290)
         );
  AOI221_X1 U2762 ( .B1(n18375), .B2(net535481), .C1(n18372), .C2(net591544), 
        .A(n4304), .ZN(n4289) );
  NAND4_X1 U2763 ( .A1(n4270), .A2(n4271), .A3(n4272), .A4(n4273), .ZN(n2774)
         );
  AOI221_X1 U2764 ( .B1(n18363), .B2(net366965), .C1(n18360), .C2(net591801), 
        .A(n4287), .ZN(n4270) );
  NOR4_X1 U2765 ( .A1(n4282), .A2(n4283), .A3(n4284), .A4(n4285), .ZN(n4272)
         );
  AOI221_X1 U2766 ( .B1(n18375), .B2(net535482), .C1(n18372), .C2(net591545), 
        .A(n4286), .ZN(n4271) );
  NAND4_X1 U2767 ( .A1(n4252), .A2(n4253), .A3(n4254), .A4(n4255), .ZN(n2775)
         );
  AOI221_X1 U2768 ( .B1(n18363), .B2(net366966), .C1(n18360), .C2(net591802), 
        .A(n4269), .ZN(n4252) );
  NOR4_X1 U2769 ( .A1(n4264), .A2(n4265), .A3(n4266), .A4(n4267), .ZN(n4254)
         );
  AOI221_X1 U2770 ( .B1(n18375), .B2(net535483), .C1(n18372), .C2(net591546), 
        .A(n4268), .ZN(n4253) );
  NAND4_X1 U2771 ( .A1(n4234), .A2(n4235), .A3(n4236), .A4(n4237), .ZN(n2776)
         );
  AOI221_X1 U2772 ( .B1(n18363), .B2(net366967), .C1(n18360), .C2(net591803), 
        .A(n4251), .ZN(n4234) );
  NOR4_X1 U2773 ( .A1(n4246), .A2(n4247), .A3(n4248), .A4(n4249), .ZN(n4236)
         );
  AOI221_X1 U2774 ( .B1(n18375), .B2(net535484), .C1(n18372), .C2(net591547), 
        .A(n4250), .ZN(n4235) );
  NAND4_X1 U2775 ( .A1(n4216), .A2(n4217), .A3(n4218), .A4(n4219), .ZN(n2777)
         );
  AOI221_X1 U2776 ( .B1(n18363), .B2(net366968), .C1(n18360), .C2(net591804), 
        .A(n4233), .ZN(n4216) );
  NOR4_X1 U2777 ( .A1(n4228), .A2(n4229), .A3(n4230), .A4(n4231), .ZN(n4218)
         );
  AOI221_X1 U2778 ( .B1(n18375), .B2(net535485), .C1(n18372), .C2(net591548), 
        .A(n4232), .ZN(n4217) );
  NAND4_X1 U2779 ( .A1(n4198), .A2(n4199), .A3(n4200), .A4(n4201), .ZN(n2778)
         );
  AOI221_X1 U2780 ( .B1(n18363), .B2(net366969), .C1(n18360), .C2(net591805), 
        .A(n4215), .ZN(n4198) );
  NOR4_X1 U2781 ( .A1(n4210), .A2(n4211), .A3(n4212), .A4(n4213), .ZN(n4200)
         );
  AOI221_X1 U2782 ( .B1(n18375), .B2(net535486), .C1(n18372), .C2(net591549), 
        .A(n4214), .ZN(n4199) );
  NAND4_X1 U2783 ( .A1(n4180), .A2(n4181), .A3(n4182), .A4(n4183), .ZN(n2779)
         );
  AOI221_X1 U2784 ( .B1(n18363), .B2(net366970), .C1(n18360), .C2(net591806), 
        .A(n4197), .ZN(n4180) );
  NOR4_X1 U2785 ( .A1(n4192), .A2(n4193), .A3(n4194), .A4(n4195), .ZN(n4182)
         );
  AOI221_X1 U2786 ( .B1(n18375), .B2(net535487), .C1(n18372), .C2(net591550), 
        .A(n4196), .ZN(n4181) );
  NAND4_X1 U2787 ( .A1(n4162), .A2(n4163), .A3(n4164), .A4(n4165), .ZN(n2780)
         );
  AOI221_X1 U2788 ( .B1(n18363), .B2(net366971), .C1(n18360), .C2(net591807), 
        .A(n4179), .ZN(n4162) );
  NOR4_X1 U2789 ( .A1(n4174), .A2(n4175), .A3(n4176), .A4(n4177), .ZN(n4164)
         );
  AOI221_X1 U2790 ( .B1(n18375), .B2(net535488), .C1(n18372), .C2(net591551), 
        .A(n4178), .ZN(n4163) );
  NAND4_X1 U2791 ( .A1(n4144), .A2(n4145), .A3(n4146), .A4(n4147), .ZN(n2781)
         );
  AOI221_X1 U2792 ( .B1(n18363), .B2(net366972), .C1(n18360), .C2(net591808), 
        .A(n4161), .ZN(n4144) );
  NOR4_X1 U2793 ( .A1(n4156), .A2(n4157), .A3(n4158), .A4(n4159), .ZN(n4146)
         );
  AOI221_X1 U2794 ( .B1(n18375), .B2(net535489), .C1(n18372), .C2(net591552), 
        .A(n4160), .ZN(n4145) );
  NAND4_X1 U2795 ( .A1(n4126), .A2(n4127), .A3(n4128), .A4(n4129), .ZN(n2782)
         );
  AOI221_X1 U2796 ( .B1(n18363), .B2(net366973), .C1(n18360), .C2(net591809), 
        .A(n4143), .ZN(n4126) );
  NOR4_X1 U2797 ( .A1(n4138), .A2(n4139), .A3(n4140), .A4(n4141), .ZN(n4128)
         );
  AOI221_X1 U2798 ( .B1(n18375), .B2(net535490), .C1(n18372), .C2(net591553), 
        .A(n4142), .ZN(n4127) );
  NAND4_X1 U2799 ( .A1(n4108), .A2(n4109), .A3(n4110), .A4(n4111), .ZN(n2783)
         );
  AOI221_X1 U2800 ( .B1(n18363), .B2(net366974), .C1(n18360), .C2(net591810), 
        .A(n4125), .ZN(n4108) );
  NOR4_X1 U2801 ( .A1(n4120), .A2(n4121), .A3(n4122), .A4(n4123), .ZN(n4110)
         );
  AOI221_X1 U2802 ( .B1(n18375), .B2(net535491), .C1(n18372), .C2(net591554), 
        .A(n4124), .ZN(n4109) );
  NAND4_X1 U2803 ( .A1(n4090), .A2(n4091), .A3(n4092), .A4(n4093), .ZN(n2784)
         );
  AOI221_X1 U2804 ( .B1(n18364), .B2(net366975), .C1(n18361), .C2(net591811), 
        .A(n4107), .ZN(n4090) );
  NOR4_X1 U2805 ( .A1(n4102), .A2(n4103), .A3(n4104), .A4(n4105), .ZN(n4092)
         );
  AOI221_X1 U2806 ( .B1(n18376), .B2(net535492), .C1(n18373), .C2(net591555), 
        .A(n4106), .ZN(n4091) );
  NAND4_X1 U2807 ( .A1(n4072), .A2(n4073), .A3(n4074), .A4(n4075), .ZN(n2785)
         );
  AOI221_X1 U2808 ( .B1(n18364), .B2(net366976), .C1(n18361), .C2(net591812), 
        .A(n4089), .ZN(n4072) );
  NOR4_X1 U2809 ( .A1(n4084), .A2(n4085), .A3(n4086), .A4(n4087), .ZN(n4074)
         );
  AOI221_X1 U2810 ( .B1(n18376), .B2(net535493), .C1(n18373), .C2(net591556), 
        .A(n4088), .ZN(n4073) );
  NAND4_X1 U2811 ( .A1(n4054), .A2(n4055), .A3(n4056), .A4(n4057), .ZN(n2786)
         );
  AOI221_X1 U2812 ( .B1(n18364), .B2(net366977), .C1(n18361), .C2(net591813), 
        .A(n4071), .ZN(n4054) );
  NOR4_X1 U2813 ( .A1(n4066), .A2(n4067), .A3(n4068), .A4(n4069), .ZN(n4056)
         );
  AOI221_X1 U2814 ( .B1(n18376), .B2(net535494), .C1(n18373), .C2(net591557), 
        .A(n4070), .ZN(n4055) );
  NAND4_X1 U2815 ( .A1(n4036), .A2(n4037), .A3(n4038), .A4(n4039), .ZN(n2787)
         );
  AOI221_X1 U2816 ( .B1(n18364), .B2(net366978), .C1(n18361), .C2(net591814), 
        .A(n4053), .ZN(n4036) );
  NOR4_X1 U2817 ( .A1(n4048), .A2(n4049), .A3(n4050), .A4(n4051), .ZN(n4038)
         );
  AOI221_X1 U2818 ( .B1(n18376), .B2(net535495), .C1(n18373), .C2(net591558), 
        .A(n4052), .ZN(n4037) );
  NAND4_X1 U2819 ( .A1(n4018), .A2(n4019), .A3(n4020), .A4(n4021), .ZN(n2788)
         );
  AOI221_X1 U2820 ( .B1(n18364), .B2(net366979), .C1(n18361), .C2(net591815), 
        .A(n4035), .ZN(n4018) );
  NOR4_X1 U2821 ( .A1(n4030), .A2(n4031), .A3(n4032), .A4(n4033), .ZN(n4020)
         );
  AOI221_X1 U2822 ( .B1(n18376), .B2(net535496), .C1(n18373), .C2(net591559), 
        .A(n4034), .ZN(n4019) );
  NAND4_X1 U2823 ( .A1(n4000), .A2(n4001), .A3(n4002), .A4(n4003), .ZN(n2789)
         );
  AOI221_X1 U2824 ( .B1(n18364), .B2(net366980), .C1(n18361), .C2(net591816), 
        .A(n4017), .ZN(n4000) );
  NOR4_X1 U2825 ( .A1(n4012), .A2(n4013), .A3(n4014), .A4(n4015), .ZN(n4002)
         );
  AOI221_X1 U2826 ( .B1(n18376), .B2(net535497), .C1(n18373), .C2(net591560), 
        .A(n4016), .ZN(n4001) );
  NAND4_X1 U2827 ( .A1(n3982), .A2(n3983), .A3(n3984), .A4(n3985), .ZN(n2790)
         );
  AOI221_X1 U2828 ( .B1(n18364), .B2(net366981), .C1(n18361), .C2(net591817), 
        .A(n3999), .ZN(n3982) );
  NOR4_X1 U2829 ( .A1(n3994), .A2(n3995), .A3(n3996), .A4(n3997), .ZN(n3984)
         );
  AOI221_X1 U2830 ( .B1(n18376), .B2(net535498), .C1(n18373), .C2(net591561), 
        .A(n3998), .ZN(n3983) );
  NAND4_X1 U2831 ( .A1(n3931), .A2(n3932), .A3(n3933), .A4(n3934), .ZN(n2791)
         );
  AOI221_X1 U2832 ( .B1(n18364), .B2(net366982), .C1(n18361), .C2(net591818), 
        .A(n3979), .ZN(n3931) );
  NOR4_X1 U2833 ( .A1(n3959), .A2(n3960), .A3(n3961), .A4(n3962), .ZN(n3933)
         );
  AOI221_X1 U2834 ( .B1(n18376), .B2(net535499), .C1(n18373), .C2(net591562), 
        .A(n3974), .ZN(n3932) );
  NAND4_X1 U2835 ( .A1(n3896), .A2(n3897), .A3(n3898), .A4(n3899), .ZN(n2792)
         );
  AOI221_X1 U2836 ( .B1(n18472), .B2(net479345), .C1(n18469), .C2(net535532), 
        .A(n3927), .ZN(n3897) );
  AOI221_X1 U2837 ( .B1(n18460), .B2(net310470), .C1(n18457), .C2(net423334), 
        .A(n3930), .ZN(n3896) );
  NOR4_X1 U2838 ( .A1(n3920), .A2(n3921), .A3(n3922), .A4(n3923), .ZN(n3898)
         );
  NAND4_X1 U2839 ( .A1(n3877), .A2(n3878), .A3(n3879), .A4(n3880), .ZN(n2794)
         );
  AOI221_X1 U2840 ( .B1(n18472), .B2(net479346), .C1(n18469), .C2(net535533), 
        .A(n3893), .ZN(n3878) );
  AOI221_X1 U2841 ( .B1(n18460), .B2(net310471), .C1(n18457), .C2(net423335), 
        .A(n3894), .ZN(n3877) );
  NOR4_X1 U2842 ( .A1(n3889), .A2(n3890), .A3(n3891), .A4(n3892), .ZN(n3879)
         );
  NAND4_X1 U2843 ( .A1(n3858), .A2(n3859), .A3(n3860), .A4(n3861), .ZN(n2796)
         );
  AOI221_X1 U2844 ( .B1(n18472), .B2(net479347), .C1(n18469), .C2(net535534), 
        .A(n3874), .ZN(n3859) );
  AOI221_X1 U2845 ( .B1(n18460), .B2(net310472), .C1(n18457), .C2(net423336), 
        .A(n3875), .ZN(n3858) );
  NOR4_X1 U2846 ( .A1(n3870), .A2(n3871), .A3(n3872), .A4(n3873), .ZN(n3860)
         );
  NAND4_X1 U2847 ( .A1(n2751), .A2(n2752), .A3(n2753), .A4(n2754), .ZN(n2798)
         );
  AOI221_X1 U2848 ( .B1(n18472), .B2(net479348), .C1(n18469), .C2(net535535), 
        .A(n3855), .ZN(n2752) );
  AOI221_X1 U2849 ( .B1(n18460), .B2(net310473), .C1(n18457), .C2(net423337), 
        .A(n3856), .ZN(n2751) );
  NOR4_X1 U2850 ( .A1(n3851), .A2(n3852), .A3(n3853), .A4(n3854), .ZN(n2753)
         );
  NAND4_X1 U2851 ( .A1(n2732), .A2(n2733), .A3(n2734), .A4(n2735), .ZN(n2800)
         );
  AOI221_X1 U2852 ( .B1(n18472), .B2(net479349), .C1(n18469), .C2(net535536), 
        .A(n2748), .ZN(n2733) );
  AOI221_X1 U2853 ( .B1(n18460), .B2(net310474), .C1(n18457), .C2(net423338), 
        .A(n2749), .ZN(n2732) );
  NOR4_X1 U2854 ( .A1(n2744), .A2(n2745), .A3(n2746), .A4(n2747), .ZN(n2734)
         );
  NAND4_X1 U2855 ( .A1(n2713), .A2(n2714), .A3(n2715), .A4(n2716), .ZN(n2802)
         );
  AOI221_X1 U2856 ( .B1(n18472), .B2(net479350), .C1(n18469), .C2(net535537), 
        .A(n2729), .ZN(n2714) );
  AOI221_X1 U2857 ( .B1(n18460), .B2(net310475), .C1(n18457), .C2(net423339), 
        .A(n2730), .ZN(n2713) );
  NOR4_X1 U2858 ( .A1(n2725), .A2(n2726), .A3(n2727), .A4(n2728), .ZN(n2715)
         );
  NAND4_X1 U2859 ( .A1(n2694), .A2(n2695), .A3(n2696), .A4(n2697), .ZN(n2804)
         );
  AOI221_X1 U2860 ( .B1(n18472), .B2(net479351), .C1(n18469), .C2(net535538), 
        .A(n2710), .ZN(n2695) );
  AOI221_X1 U2861 ( .B1(n18460), .B2(net310476), .C1(n18457), .C2(net423340), 
        .A(n2711), .ZN(n2694) );
  NOR4_X1 U2862 ( .A1(n2706), .A2(n2707), .A3(n2708), .A4(n2709), .ZN(n2696)
         );
  NAND4_X1 U2863 ( .A1(n2675), .A2(n2676), .A3(n2677), .A4(n2678), .ZN(n2806)
         );
  AOI221_X1 U2864 ( .B1(n18472), .B2(net479352), .C1(n18469), .C2(net535539), 
        .A(n2691), .ZN(n2676) );
  AOI221_X1 U2865 ( .B1(n18460), .B2(net310477), .C1(n18457), .C2(net423341), 
        .A(n2692), .ZN(n2675) );
  NOR4_X1 U2866 ( .A1(n2687), .A2(n2688), .A3(n2689), .A4(n2690), .ZN(n2677)
         );
  NAND4_X1 U2867 ( .A1(n2656), .A2(n2657), .A3(n2658), .A4(n2659), .ZN(n2808)
         );
  AOI221_X1 U2868 ( .B1(n18472), .B2(net479353), .C1(n18469), .C2(net535540), 
        .A(n2672), .ZN(n2657) );
  AOI221_X1 U2869 ( .B1(n18460), .B2(net310478), .C1(n18457), .C2(net423342), 
        .A(n2673), .ZN(n2656) );
  NOR4_X1 U2870 ( .A1(n2668), .A2(n2669), .A3(n2670), .A4(n2671), .ZN(n2658)
         );
  NAND4_X1 U2871 ( .A1(n2637), .A2(n2638), .A3(n2639), .A4(n2640), .ZN(n2810)
         );
  AOI221_X1 U2872 ( .B1(n18472), .B2(net479354), .C1(n18469), .C2(net535541), 
        .A(n2653), .ZN(n2638) );
  AOI221_X1 U2873 ( .B1(n18460), .B2(net310479), .C1(n18457), .C2(net423343), 
        .A(n2654), .ZN(n2637) );
  NOR4_X1 U2874 ( .A1(n2649), .A2(n2650), .A3(n2651), .A4(n2652), .ZN(n2639)
         );
  NAND4_X1 U2875 ( .A1(n2618), .A2(n2619), .A3(n2620), .A4(n2621), .ZN(n2812)
         );
  AOI221_X1 U2876 ( .B1(n18472), .B2(net479355), .C1(n18469), .C2(net535542), 
        .A(n2634), .ZN(n2619) );
  AOI221_X1 U2877 ( .B1(n18460), .B2(net310480), .C1(n18457), .C2(net423344), 
        .A(n2635), .ZN(n2618) );
  NOR4_X1 U2878 ( .A1(n2630), .A2(n2631), .A3(n2632), .A4(n2633), .ZN(n2620)
         );
  NAND4_X1 U2879 ( .A1(n2599), .A2(n2600), .A3(n2601), .A4(n2602), .ZN(n2814)
         );
  AOI221_X1 U2880 ( .B1(n18472), .B2(net479356), .C1(n18469), .C2(net535543), 
        .A(n2615), .ZN(n2600) );
  AOI221_X1 U2881 ( .B1(n18460), .B2(net310481), .C1(n18457), .C2(net423345), 
        .A(n2616), .ZN(n2599) );
  NOR4_X1 U2882 ( .A1(n2611), .A2(n2612), .A3(n2613), .A4(n2614), .ZN(n2601)
         );
  NAND4_X1 U2883 ( .A1(n2580), .A2(n2581), .A3(n2582), .A4(n2583), .ZN(n2816)
         );
  AOI221_X1 U2884 ( .B1(n18473), .B2(net479357), .C1(n18470), .C2(net535544), 
        .A(n2596), .ZN(n2581) );
  AOI221_X1 U2885 ( .B1(n18461), .B2(net310482), .C1(n18458), .C2(net423346), 
        .A(n2597), .ZN(n2580) );
  NOR4_X1 U2886 ( .A1(n2592), .A2(n2593), .A3(n2594), .A4(n2595), .ZN(n2582)
         );
  NAND4_X1 U2887 ( .A1(n2561), .A2(n2562), .A3(n2563), .A4(n2564), .ZN(n2818)
         );
  AOI221_X1 U2888 ( .B1(n18473), .B2(net479358), .C1(n18470), .C2(net535545), 
        .A(n2577), .ZN(n2562) );
  AOI221_X1 U2889 ( .B1(n18461), .B2(net310483), .C1(n18458), .C2(net423347), 
        .A(n2578), .ZN(n2561) );
  NOR4_X1 U2890 ( .A1(n2573), .A2(n2574), .A3(n2575), .A4(n2576), .ZN(n2563)
         );
  NAND4_X1 U2891 ( .A1(n2542), .A2(n2543), .A3(n2544), .A4(n2545), .ZN(n2820)
         );
  AOI221_X1 U2892 ( .B1(n18473), .B2(net479359), .C1(n18470), .C2(net535546), 
        .A(n2558), .ZN(n2543) );
  AOI221_X1 U2893 ( .B1(n18461), .B2(net310484), .C1(n18458), .C2(net423348), 
        .A(n2559), .ZN(n2542) );
  NOR4_X1 U2894 ( .A1(n2554), .A2(n2555), .A3(n2556), .A4(n2557), .ZN(n2544)
         );
  NAND4_X1 U2895 ( .A1(n2523), .A2(n2524), .A3(n2525), .A4(n2526), .ZN(n2822)
         );
  AOI221_X1 U2896 ( .B1(n18473), .B2(net479360), .C1(n18470), .C2(net535547), 
        .A(n2539), .ZN(n2524) );
  AOI221_X1 U2897 ( .B1(n18461), .B2(net310485), .C1(n18458), .C2(net423349), 
        .A(n2540), .ZN(n2523) );
  NOR4_X1 U2898 ( .A1(n2535), .A2(n2536), .A3(n2537), .A4(n2538), .ZN(n2525)
         );
  NAND4_X1 U2899 ( .A1(n2504), .A2(n2505), .A3(n2506), .A4(n2507), .ZN(n2824)
         );
  AOI221_X1 U2900 ( .B1(n18473), .B2(net479361), .C1(n18470), .C2(net535548), 
        .A(n2520), .ZN(n2505) );
  AOI221_X1 U2901 ( .B1(n18461), .B2(net310486), .C1(n18458), .C2(net423350), 
        .A(n2521), .ZN(n2504) );
  NOR4_X1 U2902 ( .A1(n2516), .A2(n2517), .A3(n2518), .A4(n2519), .ZN(n2506)
         );
  NAND4_X1 U2903 ( .A1(n2485), .A2(n2486), .A3(n2487), .A4(n2488), .ZN(n2826)
         );
  AOI221_X1 U2904 ( .B1(n18473), .B2(net479362), .C1(n18470), .C2(net535549), 
        .A(n2501), .ZN(n2486) );
  AOI221_X1 U2905 ( .B1(n18461), .B2(net310487), .C1(n18458), .C2(net423351), 
        .A(n2502), .ZN(n2485) );
  NOR4_X1 U2906 ( .A1(n2497), .A2(n2498), .A3(n2499), .A4(n2500), .ZN(n2487)
         );
  NAND4_X1 U2907 ( .A1(n2466), .A2(n2467), .A3(n2468), .A4(n2469), .ZN(n2828)
         );
  AOI221_X1 U2908 ( .B1(n18473), .B2(net479363), .C1(n18470), .C2(net535550), 
        .A(n2482), .ZN(n2467) );
  AOI221_X1 U2909 ( .B1(n18461), .B2(net310488), .C1(n18458), .C2(net423352), 
        .A(n2483), .ZN(n2466) );
  NOR4_X1 U2910 ( .A1(n2478), .A2(n2479), .A3(n2480), .A4(n2481), .ZN(n2468)
         );
  NAND4_X1 U2911 ( .A1(n2447), .A2(n2448), .A3(n2449), .A4(n2450), .ZN(n2830)
         );
  AOI221_X1 U2912 ( .B1(n18473), .B2(net479364), .C1(n18470), .C2(net535551), 
        .A(n2463), .ZN(n2448) );
  AOI221_X1 U2913 ( .B1(n18461), .B2(net310489), .C1(n18458), .C2(net423353), 
        .A(n2464), .ZN(n2447) );
  NOR4_X1 U2914 ( .A1(n2459), .A2(n2460), .A3(n2461), .A4(n2462), .ZN(n2449)
         );
  NAND4_X1 U2915 ( .A1(n2428), .A2(n2429), .A3(n2430), .A4(n2431), .ZN(n2832)
         );
  AOI221_X1 U2916 ( .B1(n18473), .B2(net479365), .C1(n18470), .C2(net535552), 
        .A(n2444), .ZN(n2429) );
  AOI221_X1 U2917 ( .B1(n18461), .B2(net310490), .C1(n18458), .C2(net423354), 
        .A(n2445), .ZN(n2428) );
  NOR4_X1 U2918 ( .A1(n2440), .A2(n2441), .A3(n2442), .A4(n2443), .ZN(n2430)
         );
  NAND4_X1 U2919 ( .A1(n2409), .A2(n2410), .A3(n2411), .A4(n2412), .ZN(n2834)
         );
  AOI221_X1 U2920 ( .B1(n18473), .B2(net479366), .C1(n18470), .C2(net535553), 
        .A(n2425), .ZN(n2410) );
  AOI221_X1 U2921 ( .B1(n18461), .B2(net310491), .C1(n18458), .C2(net423355), 
        .A(n2426), .ZN(n2409) );
  NOR4_X1 U2922 ( .A1(n2421), .A2(n2422), .A3(n2423), .A4(n2424), .ZN(n2411)
         );
  NAND4_X1 U2923 ( .A1(n2390), .A2(n2391), .A3(n2392), .A4(n2393), .ZN(n2836)
         );
  AOI221_X1 U2924 ( .B1(n18473), .B2(net479367), .C1(n18470), .C2(net535554), 
        .A(n2406), .ZN(n2391) );
  AOI221_X1 U2925 ( .B1(n18461), .B2(net310492), .C1(n18458), .C2(net423356), 
        .A(n2407), .ZN(n2390) );
  NOR4_X1 U2926 ( .A1(n2402), .A2(n2403), .A3(n2404), .A4(n2405), .ZN(n2392)
         );
  NAND4_X1 U2927 ( .A1(n2371), .A2(n2372), .A3(n2373), .A4(n2374), .ZN(n2838)
         );
  AOI221_X1 U2928 ( .B1(n18473), .B2(net479368), .C1(n18470), .C2(net535555), 
        .A(n2387), .ZN(n2372) );
  AOI221_X1 U2929 ( .B1(n18461), .B2(net310493), .C1(n18458), .C2(net423357), 
        .A(n2388), .ZN(n2371) );
  NOR4_X1 U2930 ( .A1(n2383), .A2(n2384), .A3(n2385), .A4(n2386), .ZN(n2373)
         );
  NAND4_X1 U2931 ( .A1(n2352), .A2(n2353), .A3(n2354), .A4(n2355), .ZN(n2840)
         );
  AOI221_X1 U2932 ( .B1(n18474), .B2(net479369), .C1(n18471), .C2(net535556), 
        .A(n2368), .ZN(n2353) );
  AOI221_X1 U2933 ( .B1(n18462), .B2(net310494), .C1(n18459), .C2(net423358), 
        .A(n2369), .ZN(n2352) );
  NOR4_X1 U2934 ( .A1(n2364), .A2(n2365), .A3(n2366), .A4(n2367), .ZN(n2354)
         );
  NAND4_X1 U2935 ( .A1(n2333), .A2(n2334), .A3(n2335), .A4(n2336), .ZN(n2842)
         );
  AOI221_X1 U2936 ( .B1(n18474), .B2(net479370), .C1(n18471), .C2(net535557), 
        .A(n2349), .ZN(n2334) );
  AOI221_X1 U2937 ( .B1(n18462), .B2(net310495), .C1(n18459), .C2(net423359), 
        .A(n2350), .ZN(n2333) );
  NOR4_X1 U2938 ( .A1(n2345), .A2(n2346), .A3(n2347), .A4(n2348), .ZN(n2335)
         );
  NAND4_X1 U2939 ( .A1(n2314), .A2(n2315), .A3(n2316), .A4(n2317), .ZN(n2844)
         );
  AOI221_X1 U2940 ( .B1(n18474), .B2(net479371), .C1(n18471), .C2(net535558), 
        .A(n2330), .ZN(n2315) );
  AOI221_X1 U2941 ( .B1(n18462), .B2(net310496), .C1(n18459), .C2(net423360), 
        .A(n2331), .ZN(n2314) );
  NOR4_X1 U2942 ( .A1(n2326), .A2(n2327), .A3(n2328), .A4(n2329), .ZN(n2316)
         );
  NAND4_X1 U2943 ( .A1(n2295), .A2(n2296), .A3(n2297), .A4(n2298), .ZN(n2846)
         );
  AOI221_X1 U2944 ( .B1(n18474), .B2(net479372), .C1(n18471), .C2(net535559), 
        .A(n2311), .ZN(n2296) );
  AOI221_X1 U2945 ( .B1(n18462), .B2(net310497), .C1(n18459), .C2(net423361), 
        .A(n2312), .ZN(n2295) );
  NOR4_X1 U2946 ( .A1(n2307), .A2(n2308), .A3(n2309), .A4(n2310), .ZN(n2297)
         );
  NAND4_X1 U2947 ( .A1(n2276), .A2(n2277), .A3(n2278), .A4(n2279), .ZN(n2848)
         );
  AOI221_X1 U2948 ( .B1(n18474), .B2(net479373), .C1(n18471), .C2(net535560), 
        .A(n2292), .ZN(n2277) );
  AOI221_X1 U2949 ( .B1(n18462), .B2(net310498), .C1(n18459), .C2(net423362), 
        .A(n2293), .ZN(n2276) );
  NOR4_X1 U2950 ( .A1(n2288), .A2(n2289), .A3(n2290), .A4(n2291), .ZN(n2278)
         );
  NAND4_X1 U2951 ( .A1(n2257), .A2(n2258), .A3(n2259), .A4(n2260), .ZN(n2850)
         );
  AOI221_X1 U2952 ( .B1(n18474), .B2(net479374), .C1(n18471), .C2(net535561), 
        .A(n2273), .ZN(n2258) );
  AOI221_X1 U2953 ( .B1(n18462), .B2(net310499), .C1(n18459), .C2(net423363), 
        .A(n2274), .ZN(n2257) );
  NOR4_X1 U2954 ( .A1(n2269), .A2(n2270), .A3(n2271), .A4(n2272), .ZN(n2259)
         );
  NAND4_X1 U2955 ( .A1(n2238), .A2(n2239), .A3(n2240), .A4(n2241), .ZN(n2852)
         );
  AOI221_X1 U2956 ( .B1(n18474), .B2(net479375), .C1(n18471), .C2(net535562), 
        .A(n2254), .ZN(n2239) );
  AOI221_X1 U2957 ( .B1(n18462), .B2(net310500), .C1(n18459), .C2(net423364), 
        .A(n2255), .ZN(n2238) );
  NOR4_X1 U2958 ( .A1(n2250), .A2(n2251), .A3(n2252), .A4(n2253), .ZN(n2240)
         );
  NAND4_X1 U2959 ( .A1(n2186), .A2(n2187), .A3(n2188), .A4(n2189), .ZN(n2854)
         );
  AOI221_X1 U2960 ( .B1(n18474), .B2(net479376), .C1(n18471), .C2(net535563), 
        .A(n2229), .ZN(n2187) );
  AOI221_X1 U2961 ( .B1(n18462), .B2(net479344), .C1(n18459), .C2(net423365), 
        .A(n2234), .ZN(n2186) );
  NOR4_X1 U2962 ( .A1(n2214), .A2(n2215), .A3(n2216), .A4(n2217), .ZN(n2188)
         );
  AND3_X1 U2963 ( .A1(ENABLE), .A2(n18999), .A3(RD1), .ZN(n18352) );
  OAI22_X1 U2964 ( .A1(n18684), .A2(n18962), .B1(n1805), .B2(n18288), .ZN(
        n3200) );
  OAI22_X1 U2965 ( .A1(n18684), .A2(n18965), .B1(n18681), .B2(n18289), .ZN(
        n3201) );
  OAI22_X1 U2966 ( .A1(n18683), .A2(n18968), .B1(n18681), .B2(n18290), .ZN(
        n3202) );
  OAI22_X1 U2967 ( .A1(n18683), .A2(n18971), .B1(n18681), .B2(n18291), .ZN(
        n3203) );
  OAI22_X1 U2968 ( .A1(n18683), .A2(n18974), .B1(n18681), .B2(n18292), .ZN(
        n3204) );
  OAI22_X1 U2969 ( .A1(n18682), .A2(n18977), .B1(n18681), .B2(n18293), .ZN(
        n3205) );
  OAI22_X1 U2970 ( .A1(n18683), .A2(n18980), .B1(n18681), .B2(n18294), .ZN(
        n3206) );
  OAI22_X1 U2971 ( .A1(n18686), .A2(n18992), .B1(n1805), .B2(n18295), .ZN(
        n3207) );
  OAI22_X1 U2972 ( .A1(n18682), .A2(n1136), .B1(n18681), .B2(n18296), .ZN(
        n3176) );
  OAI22_X1 U2973 ( .A1(n18689), .A2(n1134), .B1(n18681), .B2(n18297), .ZN(
        n3177) );
  OAI22_X1 U2974 ( .A1(n18689), .A2(n1130), .B1(n18681), .B2(n18298), .ZN(
        n3179) );
  OAI22_X1 U2975 ( .A1(n18552), .A2(n18321), .B1(n18550), .B2(n18966), .ZN(
        n2843) );
  OAI22_X1 U2976 ( .A1(n18552), .A2(n18322), .B1(n18549), .B2(n18969), .ZN(
        n2845) );
  OAI22_X1 U2977 ( .A1(n18551), .A2(n18323), .B1(n18550), .B2(n18972), .ZN(
        n2847) );
  OAI22_X1 U2978 ( .A1(n18551), .A2(n18324), .B1(n18549), .B2(n18975), .ZN(
        n2849) );
  OAI22_X1 U2979 ( .A1(n18551), .A2(n18325), .B1(n18550), .B2(n18978), .ZN(
        n2851) );
  OAI22_X1 U2980 ( .A1(n18551), .A2(n18326), .B1(n18549), .B2(n18981), .ZN(
        n2853) );
  OAI22_X1 U2981 ( .A1(n18551), .A2(n18320), .B1(n18549), .B2(n18993), .ZN(
        n2855) );
  OAI22_X1 U2982 ( .A1(n18554), .A2(n18327), .B1(n18550), .B2(n18927), .ZN(
        n2817) );
  OAI22_X1 U2983 ( .A1(n18554), .A2(n18328), .B1(n18550), .B2(n18930), .ZN(
        n2819) );
  OAI22_X1 U2984 ( .A1(n18554), .A2(n18329), .B1(n18550), .B2(n18933), .ZN(
        n2821) );
  OAI22_X1 U2985 ( .A1(n18554), .A2(n18330), .B1(n18550), .B2(n18936), .ZN(
        n2823) );
  OAI22_X1 U2986 ( .A1(n18554), .A2(n18331), .B1(n18550), .B2(n18939), .ZN(
        n2825) );
  OAI22_X1 U2987 ( .A1(n18553), .A2(n18332), .B1(n18550), .B2(n18942), .ZN(
        n2827) );
  OAI22_X1 U2988 ( .A1(n18553), .A2(n18333), .B1(n18550), .B2(n18945), .ZN(
        n2829) );
  OAI22_X1 U2989 ( .A1(n18553), .A2(n18334), .B1(n18550), .B2(n18948), .ZN(
        n2831) );
  OAI22_X1 U2990 ( .A1(n18553), .A2(n18335), .B1(n18550), .B2(n18951), .ZN(
        n2833) );
  OAI22_X1 U2991 ( .A1(n18553), .A2(n18336), .B1(n18550), .B2(n18954), .ZN(
        n2835) );
  OAI22_X1 U2992 ( .A1(n18552), .A2(n18337), .B1(n18550), .B2(n18957), .ZN(
        n2837) );
  OAI22_X1 U2993 ( .A1(n18552), .A2(n18338), .B1(n18550), .B2(n18960), .ZN(
        n2839) );
  OAI22_X1 U2994 ( .A1(n18552), .A2(n18339), .B1(n18550), .B2(n18963), .ZN(
        n2841) );
  OAI22_X1 U2995 ( .A1(n18556), .A2(n18340), .B1(n18549), .B2(n18906), .ZN(
        n2803) );
  OAI22_X1 U2996 ( .A1(n18556), .A2(n18341), .B1(n18549), .B2(n18909), .ZN(
        n2805) );
  OAI22_X1 U2997 ( .A1(n18555), .A2(n18342), .B1(n18549), .B2(n18912), .ZN(
        n2807) );
  OAI22_X1 U2998 ( .A1(n18555), .A2(n18343), .B1(n18549), .B2(n18915), .ZN(
        n2809) );
  OAI22_X1 U2999 ( .A1(n18555), .A2(n18344), .B1(n18549), .B2(n18918), .ZN(
        n2811) );
  OAI22_X1 U3000 ( .A1(n18555), .A2(n18345), .B1(n18549), .B2(n18921), .ZN(
        n2813) );
  OAI22_X1 U3001 ( .A1(n18555), .A2(n18346), .B1(n18549), .B2(n18924), .ZN(
        n2815) );
  OAI22_X1 U3002 ( .A1(n1282), .A2(n18682), .B1(n18681), .B2(n18299), .ZN(
        n3178) );
  OAI22_X1 U3003 ( .A1(n1694), .A2(n18682), .B1(n18681), .B2(n18300), .ZN(
        n3180) );
  OAI22_X1 U3004 ( .A1(n18689), .A2(n18905), .B1(n18681), .B2(n18301), .ZN(
        n3181) );
  OAI22_X1 U3005 ( .A1(n18689), .A2(n18908), .B1(n18681), .B2(n18302), .ZN(
        n3182) );
  OAI22_X1 U3006 ( .A1(n18688), .A2(n18911), .B1(n18681), .B2(n18303), .ZN(
        n3183) );
  OAI22_X1 U3007 ( .A1(n18688), .A2(n18914), .B1(n18681), .B2(n18304), .ZN(
        n3184) );
  OAI22_X1 U3008 ( .A1(n18688), .A2(n18917), .B1(n18681), .B2(n18305), .ZN(
        n3185) );
  OAI22_X1 U3009 ( .A1(n18688), .A2(n18920), .B1(n18681), .B2(n18306), .ZN(
        n3186) );
  OAI22_X1 U3010 ( .A1(n18687), .A2(n18923), .B1(n18681), .B2(n18307), .ZN(
        n3187) );
  OAI22_X1 U3011 ( .A1(n18687), .A2(n18926), .B1(n1805), .B2(n18308), .ZN(
        n3188) );
  OAI22_X1 U3012 ( .A1(n18687), .A2(n18929), .B1(n1805), .B2(n18309), .ZN(
        n3189) );
  OAI22_X1 U3013 ( .A1(n18687), .A2(n18932), .B1(n1805), .B2(n18310), .ZN(
        n3190) );
  OAI22_X1 U3014 ( .A1(n18686), .A2(n18935), .B1(n1805), .B2(n18311), .ZN(
        n3191) );
  OAI22_X1 U3015 ( .A1(n18686), .A2(n18938), .B1(n1805), .B2(n18312), .ZN(
        n3192) );
  OAI22_X1 U3016 ( .A1(n18686), .A2(n18941), .B1(n1805), .B2(n18313), .ZN(
        n3193) );
  OAI22_X1 U3017 ( .A1(n18685), .A2(n18944), .B1(n1805), .B2(n18314), .ZN(
        n3194) );
  OAI22_X1 U3018 ( .A1(n18685), .A2(n18947), .B1(n1805), .B2(n18315), .ZN(
        n3195) );
  OAI22_X1 U3019 ( .A1(n18685), .A2(n18950), .B1(n1805), .B2(n18316), .ZN(
        n3196) );
  OAI22_X1 U3020 ( .A1(n18685), .A2(n18953), .B1(n18681), .B2(n18317), .ZN(
        n3197) );
  OAI22_X1 U3021 ( .A1(n18684), .A2(n18956), .B1(n18681), .B2(n18318), .ZN(
        n3198) );
  OAI22_X1 U3022 ( .A1(n18684), .A2(n18959), .B1(n18681), .B2(n18319), .ZN(
        n3199) );
  OAI22_X1 U3023 ( .A1(n18557), .A2(n18347), .B1(n1174), .B2(n18549), .ZN(
        n2793) );
  OAI22_X1 U3024 ( .A1(n18557), .A2(n18348), .B1(n1209), .B2(n18549), .ZN(
        n2795) );
  OAI22_X1 U3025 ( .A1(n18556), .A2(n18349), .B1(n1282), .B2(n18549), .ZN(
        n2797) );
  OAI22_X1 U3026 ( .A1(n18556), .A2(n18350), .B1(n1419), .B2(n18549), .ZN(
        n2799) );
  OAI22_X1 U3027 ( .A1(n18556), .A2(n18351), .B1(n1694), .B2(n18549), .ZN(
        n2801) );
  NAND2_X1 U3028 ( .A1(DATAIN[5]), .A2(n18999), .ZN(n1126) );
  NAND2_X1 U3029 ( .A1(DATAIN[6]), .A2(n18997), .ZN(n1124) );
  NAND2_X1 U3030 ( .A1(DATAIN[7]), .A2(n18999), .ZN(n1122) );
  NAND2_X1 U3031 ( .A1(DATAIN[8]), .A2(n18998), .ZN(n1120) );
  NAND2_X1 U3032 ( .A1(DATAIN[9]), .A2(n18997), .ZN(n1118) );
  NAND2_X1 U3033 ( .A1(DATAIN[10]), .A2(n18998), .ZN(n1116) );
  NAND2_X1 U3034 ( .A1(DATAIN[11]), .A2(n18999), .ZN(n1114) );
  NAND2_X1 U3035 ( .A1(DATAIN[12]), .A2(n18999), .ZN(n1112) );
  NAND2_X1 U3036 ( .A1(DATAIN[13]), .A2(n18998), .ZN(n1110) );
  NAND2_X1 U3037 ( .A1(DATAIN[14]), .A2(n18997), .ZN(n1108) );
  NAND2_X1 U3038 ( .A1(DATAIN[15]), .A2(n18997), .ZN(n1106) );
  NAND2_X1 U3039 ( .A1(DATAIN[16]), .A2(n18998), .ZN(n1104) );
  NAND2_X1 U3040 ( .A1(DATAIN[17]), .A2(n18997), .ZN(n1102) );
  NAND2_X1 U3041 ( .A1(DATAIN[18]), .A2(n18998), .ZN(n1100) );
  NAND2_X1 U3042 ( .A1(DATAIN[19]), .A2(n18998), .ZN(n1098) );
  NAND2_X1 U3043 ( .A1(DATAIN[20]), .A2(n18998), .ZN(n1096) );
  NAND2_X1 U3044 ( .A1(DATAIN[21]), .A2(n18999), .ZN(n1094) );
  NAND2_X1 U3045 ( .A1(DATAIN[22]), .A2(n18997), .ZN(n1092) );
  NAND2_X1 U3046 ( .A1(DATAIN[23]), .A2(n18997), .ZN(n1090) );
  NAND2_X1 U3047 ( .A1(DATAIN[24]), .A2(n18999), .ZN(n1088) );
  NAND2_X1 U3048 ( .A1(DATAIN[25]), .A2(n18998), .ZN(n1086) );
  NAND2_X1 U3049 ( .A1(DATAIN[26]), .A2(n18999), .ZN(n1084) );
  NAND2_X1 U3050 ( .A1(DATAIN[27]), .A2(n18998), .ZN(n1082) );
  NAND2_X1 U3051 ( .A1(DATAIN[28]), .A2(n18997), .ZN(n1080) );
  NAND2_X1 U3052 ( .A1(DATAIN[29]), .A2(n18997), .ZN(n1078) );
  NAND2_X1 U3053 ( .A1(DATAIN[30]), .A2(n18997), .ZN(n1076) );
  NAND2_X1 U3054 ( .A1(DATAIN[31]), .A2(n18997), .ZN(n1073) );
  NAND2_X1 U3055 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .ZN(n1247) );
  NAND2_X1 U3056 ( .A1(ADD_WR[1]), .A2(n2114), .ZN(n1212) );
  NAND2_X1 U3057 ( .A1(ADD_WR[0]), .A2(n2113), .ZN(n1176) );
  AND3_X1 U3058 ( .A1(WR), .A2(ENABLE), .A3(ADD_WR[4]), .ZN(n1803) );
  AND3_X1 U3059 ( .A1(ENABLE), .A2(n1664), .A3(WR), .ZN(n1250) );
  INV_X1 U3060 ( .A(ADD_WR[4]), .ZN(n1664) );
  INV_X1 U3061 ( .A(ADD_WR[3]), .ZN(n1249) );
  INV_X1 U3062 ( .A(ADD_WR[2]), .ZN(n1248) );
  INV_X1 U3063 ( .A(ADD_WR[0]), .ZN(n2114) );
  INV_X1 U3064 ( .A(ADD_WR[1]), .ZN(n2113) );
  INV_X1 U3065 ( .A(n17839), .ZN(n18441) );
  INV_X1 U3066 ( .A(n18352), .ZN(n18539) );
endmodule


module write_back_stage ( LMD_OUT, ALU_MA_OUT, MUX_SEL_WB, RF_DATA_IN );
  input [31:0] LMD_OUT;
  input [31:0] ALU_MA_OUT;
  output [31:0] RF_DATA_IN;
  input MUX_SEL_WB;


  MUX21_GENERIC_N32_1 Mux_wb ( .A(ALU_MA_OUT), .B(LMD_OUT), .SEL(MUX_SEL_WB), 
        .Y(RF_DATA_IN) );
endmodule


module mem_access_stage ( ALU_OUT, REGB_EX_OUT, DRAM_WE, LMD_LATCH_EN, DRAM_EN, 
        RST, CLK, ALU_MA_LATCH_EN, FLUSH, ALU_MA_OUT, LMD_OUT );
  input [31:0] ALU_OUT;
  input [31:0] REGB_EX_OUT;
  output [31:0] ALU_MA_OUT;
  output [31:0] LMD_OUT;
  input DRAM_WE, LMD_LATCH_EN, DRAM_EN, RST, CLK, ALU_MA_LATCH_EN, FLUSH;
  wire   sig_wr_enable, n1, sig_fd_2, sig_fd_1;
  wire   [31:0] reg_lmd_in;
  assign n1 = RST;

  DRAM_MEM_DEPTH80_D_SIZE32 DRAM_0 ( .RESET(n1), .CLK(CLK), .DATAIN(
        REGB_EX_OUT), .ENABLE(DRAM_EN), .WR_enable(sig_wr_enable), .Addr(
        ALU_OUT), .Dout(reg_lmd_in) );
  reg_generic_N32_1 reg_lmd ( .D(reg_lmd_in), .CLK(CLK), .RST(n1), .EN(
        LMD_LATCH_EN), .Q(LMD_OUT) );
  reg_generic_N32_0 reg_alu_MA ( .D(ALU_OUT), .CLK(CLK), .RST(n1), .EN(
        ALU_MA_LATCH_EN), .Q(ALU_MA_OUT) );
  FD_s_321 ff_1 ( .D(FLUSH), .CLK(CLK), .RST(n1), .EN(1'b1), .Q(sig_fd_1) );
  FD_s_320 ff_2 ( .D(sig_fd_1), .CLK(CLK), .RST(n1), .EN(1'b1), .Q(sig_fd_2)
         );
  MUX21_1 mux_dram_flush ( .A(1'b0), .B(DRAM_WE), .SEL(sig_fd_2), .Y(
        sig_wr_enable) );
endmodule


module execute_stage ( CLK, RST, NPC_EXECUTE_IN, REGA_OUT, REGB_OUT, 
        REGIMM_OUT, ALU_OPCODE, MUX_SEL_ANPC, MUX_SEL_BIMM, MUX_SEL_JAL_IMM, 
        MUX_SEL_ALU_32, MUX_SEL_ALU_1, ALU_OUTREG_EN, REGBDELAY_LATCH_EN, 
        REGALU_OUT, REGB_EX_OUT );
  input [31:0] NPC_EXECUTE_IN;
  input [31:0] REGA_OUT;
  input [31:0] REGB_OUT;
  input [31:0] REGIMM_OUT;
  input [7:0] ALU_OPCODE;
  input [2:0] MUX_SEL_ALU_32;
  input [1:0] MUX_SEL_ALU_1;
  output [31:0] REGALU_OUT;
  output [31:0] REGB_EX_OUT;
  input CLK, RST, MUX_SEL_ANPC, MUX_SEL_BIMM, MUX_SEL_JAL_IMM, ALU_OUTREG_EN,
         REGBDELAY_LATCH_EN;
  wire   sig_ne, sig_ge, sig_le, sig_ee, \sig_comparison[0] ,
         \sig_mux_imm_4[9] , \sig_mux_imm_4[8] , \sig_mux_imm_4[7] ,
         \sig_mux_imm_4[6] , \sig_mux_imm_4[5] , \sig_mux_imm_4[4] ,
         \sig_mux_imm_4[3] , \sig_mux_imm_4[31] , \sig_mux_imm_4[30] ,
         \sig_mux_imm_4[2] , \sig_mux_imm_4[29] , \sig_mux_imm_4[28] ,
         \sig_mux_imm_4[27] , \sig_mux_imm_4[26] , \sig_mux_imm_4[25] ,
         \sig_mux_imm_4[24] , \sig_mux_imm_4[23] , \sig_mux_imm_4[22] ,
         \sig_mux_imm_4[21] , \sig_mux_imm_4[20] , \sig_mux_imm_4[1] ,
         \sig_mux_imm_4[19] , \sig_mux_imm_4[18] , \sig_mux_imm_4[17] ,
         \sig_mux_imm_4[16] , \sig_mux_imm_4[15] , \sig_mux_imm_4[14] ,
         \sig_mux_imm_4[13] , \sig_mux_imm_4[12] , \sig_mux_imm_4[11] ,
         \sig_mux_imm_4[10] , \sig_mux_imm_4[0] ;
  wire   [31:0] alu_a;
  wire   [31:0] alu_b;
  wire   [31:0] sig_add;
  wire   [31:0] sig_shift;
  wire   [31:0] sig_logic;
  wire   [31:0] sig_mult;
  wire   [31:0] reg_alu_in;

  MUX21_GENERIC_N32_4 mux_a_npc ( .A(NPC_EXECUTE_IN), .B(REGA_OUT), .SEL(
        MUX_SEL_ANPC), .Y(alu_a) );
  MUX21_GENERIC_N32_3 mux_imm_4 ( .A(REGIMM_OUT), .B({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .SEL(MUX_SEL_JAL_IMM), .Y({
        \sig_mux_imm_4[31] , \sig_mux_imm_4[30] , \sig_mux_imm_4[29] , 
        \sig_mux_imm_4[28] , \sig_mux_imm_4[27] , \sig_mux_imm_4[26] , 
        \sig_mux_imm_4[25] , \sig_mux_imm_4[24] , \sig_mux_imm_4[23] , 
        \sig_mux_imm_4[22] , \sig_mux_imm_4[21] , \sig_mux_imm_4[20] , 
        \sig_mux_imm_4[19] , \sig_mux_imm_4[18] , \sig_mux_imm_4[17] , 
        \sig_mux_imm_4[16] , \sig_mux_imm_4[15] , \sig_mux_imm_4[14] , 
        \sig_mux_imm_4[13] , \sig_mux_imm_4[12] , \sig_mux_imm_4[11] , 
        \sig_mux_imm_4[10] , \sig_mux_imm_4[9] , \sig_mux_imm_4[8] , 
        \sig_mux_imm_4[7] , \sig_mux_imm_4[6] , \sig_mux_imm_4[5] , 
        \sig_mux_imm_4[4] , \sig_mux_imm_4[3] , \sig_mux_imm_4[2] , 
        \sig_mux_imm_4[1] , \sig_mux_imm_4[0] }) );
  MUX21_GENERIC_N32_2 mux_b_imm ( .A(REGB_OUT), .B({\sig_mux_imm_4[31] , 
        \sig_mux_imm_4[30] , \sig_mux_imm_4[29] , \sig_mux_imm_4[28] , 
        \sig_mux_imm_4[27] , \sig_mux_imm_4[26] , \sig_mux_imm_4[25] , 
        \sig_mux_imm_4[24] , \sig_mux_imm_4[23] , \sig_mux_imm_4[22] , 
        \sig_mux_imm_4[21] , \sig_mux_imm_4[20] , \sig_mux_imm_4[19] , 
        \sig_mux_imm_4[18] , \sig_mux_imm_4[17] , \sig_mux_imm_4[16] , 
        \sig_mux_imm_4[15] , \sig_mux_imm_4[14] , \sig_mux_imm_4[13] , 
        \sig_mux_imm_4[12] , \sig_mux_imm_4[11] , \sig_mux_imm_4[10] , 
        \sig_mux_imm_4[9] , \sig_mux_imm_4[8] , \sig_mux_imm_4[7] , 
        \sig_mux_imm_4[6] , \sig_mux_imm_4[5] , \sig_mux_imm_4[4] , 
        \sig_mux_imm_4[3] , \sig_mux_imm_4[2] , \sig_mux_imm_4[1] , 
        \sig_mux_imm_4[0] }), .SEL(MUX_SEL_BIMM), .Y(alu_b) );
  ALU_N32 Alu_exe ( .ALU_OPCODE(ALU_OPCODE), .A(alu_a), .B(alu_b), .Y_ADDER(
        sig_add), .Y_SHIFT(sig_shift), .Y_LOGIC(sig_logic), .Y_MULT(sig_mult), 
        .ne(sig_ne), .ge(sig_ge), .le(sig_le), .ee(sig_ee) );
  MUX41_1 mux_alu_comparator ( .A(sig_ne), .B(sig_ge), .C(sig_le), .D(sig_ee), 
        .SEL(MUX_SEL_ALU_1), .Y(\sig_comparison[0] ) );
  MUX51_GENERIC_N32 mux_alu_32 ( .A(sig_add), .B(sig_logic), .C(sig_shift), 
        .D({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \sig_comparison[0] }), 
        .E(sig_mult), .SEL(MUX_SEL_ALU_32), .Y(reg_alu_in) );
  reg_generic_N32_3 reg_alu ( .D(reg_alu_in), .CLK(CLK), .RST(RST), .EN(
        ALU_OUTREG_EN), .Q(REGALU_OUT) );
  reg_generic_N32_2 regB_delay ( .D(REGB_OUT), .CLK(CLK), .RST(RST), .EN(
        REGBDELAY_LATCH_EN), .Q(REGB_EX_OUT) );
endmodule


module decode_stage ( RST, CLK, SOURCE1, SOURCE2, DESTINATION, IMMEDIATE, NPC, 
        RD1_EN, RD2_EN, WR_EN_WB, RF_DATAIN, REGA_LATCH_EN, REGB_LATCH_EN, 
        REGIMM_LATCH_EN, NPC_LATCH_DEC_EN, MUX_SEL_IMM, JUMPFC, 
        MUX_SEL_JAL_ADDR_LW, REGA_OUT, REGB_OUT, REGIMM_OUT, NPC_EXECUTE_IN, 
        NPC_DECODE_OUT, FLUSH, REG_DELAY1, REG_DELAY2, REG_DELAY3, REG_DELAY4, 
        EN_IN );
  input [4:0] SOURCE1;
  input [4:0] SOURCE2;
  input [5:0] DESTINATION;
  input [25:0] IMMEDIATE;
  input [31:0] NPC;
  input [31:0] RF_DATAIN;
  input [1:0] JUMPFC;
  input [1:0] MUX_SEL_JAL_ADDR_LW;
  output [31:0] REGA_OUT;
  output [31:0] REGB_OUT;
  output [31:0] REGIMM_OUT;
  output [31:0] NPC_EXECUTE_IN;
  output [31:0] NPC_DECODE_OUT;
  output [5:0] REG_DELAY1;
  output [5:0] REG_DELAY2;
  output [5:0] REG_DELAY3;
  output [5:0] REG_DELAY4;
  input RST, CLK, RD1_EN, RD2_EN, WR_EN_WB, REGA_LATCH_EN, REGB_LATCH_EN,
         REGIMM_LATCH_EN, NPC_LATCH_DEC_EN, MUX_SEL_IMM, EN_IN;
  output FLUSH;
  wire   sig_wr_flush, eq_cond, neq_cond, n36, n37, \sig_npc[9] , \sig_npc[8] ,
         \sig_npc[7] , \sig_npc[6] , \sig_npc[5] , \sig_npc[4] , \sig_npc[3] ,
         \sig_npc[31] , \sig_npc[30] , \sig_npc[2] , \sig_npc[29] ,
         \sig_npc[28] , \sig_npc[27] , \sig_npc[26] , \sig_npc[25] ,
         \sig_npc[24] , \sig_npc[23] , \sig_npc[22] , \sig_npc[21] ,
         \sig_npc[20] , \sig_npc[1] , \sig_npc[19] , \sig_npc[18] ,
         \sig_npc[17] , \sig_npc[16] , \sig_npc[15] , \sig_npc[14] ,
         \sig_npc[13] , \sig_npc[12] , \sig_npc[11] , \sig_npc[10] ,
         \sig_npc[0] , sig_fd_4, sig_fd_3, sig_fd_2, sig_fd_1,
         \mux_imm_out[9] , \mux_imm_out[8] , \mux_imm_out[7] ,
         \mux_imm_out[6] , \mux_imm_out[5] , \mux_imm_out[4] ,
         \mux_imm_out[3] , \mux_imm_out[31] , \mux_imm_out[30] ,
         \mux_imm_out[2] , \mux_imm_out[29] , \mux_imm_out[28] ,
         \mux_imm_out[27] , \mux_imm_out[26] , \mux_imm_out[25] ,
         \mux_imm_out[24] , \mux_imm_out[23] , \mux_imm_out[22] ,
         \mux_imm_out[21] , \mux_imm_out[20] , \mux_imm_out[1] ,
         \mux_imm_out[19] , \mux_imm_out[18] , \mux_imm_out[17] ,
         \mux_imm_out[16] , \mux_imm_out[15] , \mux_imm_out[14] ,
         \mux_imm_out[13] , \mux_imm_out[12] , \mux_imm_out[11] ,
         \mux_imm_out[10] , \mux_imm_out[0] , \addJ_out[9] , \addJ_out[8] ,
         \addJ_out[7] , \addJ_out[6] , \addJ_out[5] , \addJ_out[4] ,
         \addJ_out[3] , \addJ_out[31] , \addJ_out[30] , \addJ_out[2] ,
         \addJ_out[29] , \addJ_out[28] , \addJ_out[27] , \addJ_out[26] ,
         \addJ_out[25] , \addJ_out[24] , \addJ_out[23] , \addJ_out[22] ,
         \addJ_out[21] , \addJ_out[20] , \addJ_out[1] , \addJ_out[19] ,
         \addJ_out[18] , \addJ_out[17] , \addJ_out[16] , \addJ_out[15] ,
         \addJ_out[14] , \addJ_out[13] , \addJ_out[12] , \addJ_out[11] ,
         \addJ_out[10] , \addJ_out[0] , n40, n41, n42;
  wire   [31:0] rega_in;
  wire   [31:0] regb_in;
  wire   [25:0] sig_immediate;
  wire   [4:0] sig_source2_delay1;
  wire   [5:0] add_wr_1;
  assign n37 = RST;

  register_file_N32_A5_tot_regs32 RF ( .CLK(CLK), .RESET(n42), .ENABLE(1'b1), 
        .RD1(RD1_EN), .RD2(RD2_EN), .WR(sig_wr_flush), .ADD_WR(REG_DELAY4[4:0]), .ADD_RD1(SOURCE1), .ADD_RD2(SOURCE2), .DATAIN(RF_DATAIN), .OUT1(rega_in), 
        .OUT2(regb_in) );
  reg_generic_N26 reg_imm ( .D(IMMEDIATE), .CLK(CLK), .RST(n42), .EN(EN_IN), 
        .Q({sig_immediate[25:16], n36, sig_immediate[14:0]}) );
  reg_generic_N32_8 reg_npc_in ( .D(NPC), .CLK(CLK), .RST(n42), .EN(EN_IN), 
        .Q({\sig_npc[31] , \sig_npc[30] , \sig_npc[29] , \sig_npc[28] , 
        \sig_npc[27] , \sig_npc[26] , \sig_npc[25] , \sig_npc[24] , 
        \sig_npc[23] , \sig_npc[22] , \sig_npc[21] , \sig_npc[20] , 
        \sig_npc[19] , \sig_npc[18] , \sig_npc[17] , \sig_npc[16] , 
        \sig_npc[15] , \sig_npc[14] , \sig_npc[13] , \sig_npc[12] , 
        \sig_npc[11] , \sig_npc[10] , \sig_npc[9] , \sig_npc[8] , \sig_npc[7] , 
        \sig_npc[6] , \sig_npc[5] , \sig_npc[4] , \sig_npc[3] , \sig_npc[2] , 
        \sig_npc[1] , \sig_npc[0] }) );
  reg_generic_N5 reg_source2_delay1 ( .D(SOURCE2), .CLK(CLK), .RST(n42), .EN(
        1'b1), .Q(sig_source2_delay1) );
  reg_wr_0 reg_add_wr_delay_0 ( .D(DESTINATION), .CLK(CLK), .RST(n42), .EN(
        1'b1), .Q(REG_DELAY1) );
  MUX41_GENERIC_N6 mux_wr_rf ( .A(REG_DELAY1), .B({1'b0, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1}), .C({1'b0, sig_source2_delay1}), .D({1'b1, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .SEL(MUX_SEL_JAL_ADDR_LW), .Y(add_wr_1) );
  reg_wr_3 reg_add_wr_delay_1 ( .D(add_wr_1), .CLK(CLK), .RST(n42), .EN(1'b1), 
        .Q(REG_DELAY2) );
  reg_wr_2 reg_add_wr_delay_2 ( .D(REG_DELAY2), .CLK(CLK), .RST(n42), .EN(1'b1), .Q(REG_DELAY3) );
  reg_wr_1 reg_add_wr_delay_3 ( .D(REG_DELAY3), .CLK(CLK), .RST(n42), .EN(1'b1), .Q(REG_DELAY4) );
  zero_detector_N32 zero_det ( .A(regb_in), .YE(eq_cond) );
  MUX21_GENERIC_N32_0 mux_imm_size ( .A({n41, n40, n40, n40, n40, n40, n40, 
        n40, n40, n41, n40, n40, n40, n40, n40, n40, n40, sig_immediate[14:0]}), .B({sig_immediate[25], sig_immediate[25], sig_immediate[25], 
        sig_immediate[25], sig_immediate[25], sig_immediate[25], 
        sig_immediate[25:16], n40, sig_immediate[14:0]}), .SEL(MUX_SEL_IMM), 
        .Y({\mux_imm_out[31] , \mux_imm_out[30] , \mux_imm_out[29] , 
        \mux_imm_out[28] , \mux_imm_out[27] , \mux_imm_out[26] , 
        \mux_imm_out[25] , \mux_imm_out[24] , \mux_imm_out[23] , 
        \mux_imm_out[22] , \mux_imm_out[21] , \mux_imm_out[20] , 
        \mux_imm_out[19] , \mux_imm_out[18] , \mux_imm_out[17] , 
        \mux_imm_out[16] , \mux_imm_out[15] , \mux_imm_out[14] , 
        \mux_imm_out[13] , \mux_imm_out[12] , \mux_imm_out[11] , 
        \mux_imm_out[10] , \mux_imm_out[9] , \mux_imm_out[8] , 
        \mux_imm_out[7] , \mux_imm_out[6] , \mux_imm_out[5] , \mux_imm_out[4] , 
        \mux_imm_out[3] , \mux_imm_out[2] , \mux_imm_out[1] , \mux_imm_out[0] }) );
  P4adder_N32_M4_0 Add_J ( .A({\mux_imm_out[31] , \mux_imm_out[30] , 
        \mux_imm_out[29] , \mux_imm_out[28] , \mux_imm_out[27] , 
        \mux_imm_out[26] , \mux_imm_out[25] , \mux_imm_out[24] , 
        \mux_imm_out[23] , \mux_imm_out[22] , \mux_imm_out[21] , 
        \mux_imm_out[20] , \mux_imm_out[19] , \mux_imm_out[18] , 
        \mux_imm_out[17] , \mux_imm_out[16] , \mux_imm_out[15] , 
        \mux_imm_out[14] , \mux_imm_out[13] , \mux_imm_out[12] , 
        \mux_imm_out[11] , \mux_imm_out[10] , \mux_imm_out[9] , 
        \mux_imm_out[8] , \mux_imm_out[7] , \mux_imm_out[6] , \mux_imm_out[5] , 
        \mux_imm_out[4] , \mux_imm_out[3] , \mux_imm_out[2] , \mux_imm_out[1] , 
        \mux_imm_out[0] }), .B({\sig_npc[31] , \sig_npc[30] , \sig_npc[29] , 
        \sig_npc[28] , \sig_npc[27] , \sig_npc[26] , \sig_npc[25] , 
        \sig_npc[24] , \sig_npc[23] , \sig_npc[22] , \sig_npc[21] , 
        \sig_npc[20] , \sig_npc[19] , \sig_npc[18] , \sig_npc[17] , 
        \sig_npc[16] , \sig_npc[15] , \sig_npc[14] , \sig_npc[13] , 
        \sig_npc[12] , \sig_npc[11] , \sig_npc[10] , \sig_npc[9] , 
        \sig_npc[8] , \sig_npc[7] , \sig_npc[6] , \sig_npc[5] , \sig_npc[4] , 
        \sig_npc[3] , \sig_npc[2] , \sig_npc[1] , \sig_npc[0] }), .Y({
        \addJ_out[31] , \addJ_out[30] , \addJ_out[29] , \addJ_out[28] , 
        \addJ_out[27] , \addJ_out[26] , \addJ_out[25] , \addJ_out[24] , 
        \addJ_out[23] , \addJ_out[22] , \addJ_out[21] , \addJ_out[20] , 
        \addJ_out[19] , \addJ_out[18] , \addJ_out[17] , \addJ_out[16] , 
        \addJ_out[15] , \addJ_out[14] , \addJ_out[13] , \addJ_out[12] , 
        \addJ_out[11] , \addJ_out[10] , \addJ_out[9] , \addJ_out[8] , 
        \addJ_out[7] , \addJ_out[6] , \addJ_out[5] , \addJ_out[4] , 
        \addJ_out[3] , \addJ_out[2] , \addJ_out[1] , \addJ_out[0] }), .Ci(1'b0) );
  MUX21_GENERIC_N32_5 mux_npc_selection ( .A({\addJ_out[31] , \addJ_out[30] , 
        \addJ_out[29] , \addJ_out[28] , \addJ_out[27] , \addJ_out[26] , 
        \addJ_out[25] , \addJ_out[24] , \addJ_out[23] , \addJ_out[22] , 
        \addJ_out[21] , \addJ_out[20] , \addJ_out[19] , \addJ_out[18] , 
        \addJ_out[17] , \addJ_out[16] , \addJ_out[15] , \addJ_out[14] , 
        \addJ_out[13] , \addJ_out[12] , \addJ_out[11] , \addJ_out[10] , 
        \addJ_out[9] , \addJ_out[8] , \addJ_out[7] , \addJ_out[6] , 
        \addJ_out[5] , \addJ_out[4] , \addJ_out[3] , \addJ_out[2] , 
        \addJ_out[1] , \addJ_out[0] }), .B(NPC), .SEL(FLUSH), .Y(
        NPC_DECODE_OUT) );
  MUX41_0 mux_jump_condition_res ( .A(1'b0), .B(1'b1), .C(eq_cond), .D(
        neq_cond), .SEL(JUMPFC), .Y(FLUSH) );
  reg_generic_N32_7 reg_a ( .D(rega_in), .CLK(CLK), .RST(n42), .EN(
        REGA_LATCH_EN), .Q(REGA_OUT) );
  reg_generic_N32_6 reg_b ( .D(regb_in), .CLK(CLK), .RST(n42), .EN(
        REGB_LATCH_EN), .Q(REGB_OUT) );
  reg_generic_N32_5 regimmm ( .D({n40, n40, n40, n40, n40, n40, n40, n40, n40, 
        n40, n40, n40, n40, n40, n40, n40, n40, sig_immediate[14:0]}), .CLK(
        CLK), .RST(n42), .EN(REGIMM_LATCH_EN), .Q(REGIMM_OUT) );
  reg_generic_N32_4 reg_npc ( .D({\sig_npc[31] , \sig_npc[30] , \sig_npc[29] , 
        \sig_npc[28] , \sig_npc[27] , \sig_npc[26] , \sig_npc[25] , 
        \sig_npc[24] , \sig_npc[23] , \sig_npc[22] , \sig_npc[21] , 
        \sig_npc[20] , \sig_npc[19] , \sig_npc[18] , \sig_npc[17] , 
        \sig_npc[16] , \sig_npc[15] , \sig_npc[14] , \sig_npc[13] , 
        \sig_npc[12] , \sig_npc[11] , \sig_npc[10] , \sig_npc[9] , 
        \sig_npc[8] , \sig_npc[7] , \sig_npc[6] , \sig_npc[5] , \sig_npc[4] , 
        \sig_npc[3] , \sig_npc[2] , \sig_npc[1] , \sig_npc[0] }), .CLK(CLK), 
        .RST(n42), .EN(NPC_LATCH_DEC_EN), .Q(NPC_EXECUTE_IN) );
  FD_s_325 ff_1 ( .D(FLUSH), .CLK(CLK), .RST(n42), .EN(1'b1), .Q(sig_fd_1) );
  FD_s_324 ff_2 ( .D(sig_fd_1), .CLK(CLK), .RST(n42), .EN(1'b1), .Q(sig_fd_2)
         );
  FD_s_323 ff_3 ( .D(sig_fd_2), .CLK(CLK), .RST(n42), .EN(1'b1), .Q(sig_fd_3)
         );
  FD_s_322 ff_4 ( .D(sig_fd_3), .CLK(CLK), .RST(n42), .EN(1'b1), .Q(sig_fd_4)
         );
  MUX21_0 mux_rf_flush ( .A(1'b0), .B(WR_EN_WB), .SEL(sig_fd_4), .Y(
        sig_wr_flush) );
  INV_X1 U3 ( .A(eq_cond), .ZN(neq_cond) );
  BUF_X1 U4 ( .A(n37), .Z(n42) );
  BUF_X1 U5 ( .A(n36), .Z(n40) );
  BUF_X1 U6 ( .A(n36), .Z(n41) );
endmodule


module Add4_N32_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , n1;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];
  assign \carry[3]  = A[2];

  XOR2_X1 U3 ( .A(A[30]), .B(\carry[30] ), .Z(SUM[30]) );
  XOR2_X1 U5 ( .A(A[29]), .B(\carry[29] ), .Z(SUM[29]) );
  XOR2_X1 U7 ( .A(A[28]), .B(\carry[28] ), .Z(SUM[28]) );
  XOR2_X1 U9 ( .A(A[27]), .B(\carry[27] ), .Z(SUM[27]) );
  XOR2_X1 U11 ( .A(A[26]), .B(\carry[26] ), .Z(SUM[26]) );
  XOR2_X1 U13 ( .A(A[25]), .B(\carry[25] ), .Z(SUM[25]) );
  XOR2_X1 U15 ( .A(A[24]), .B(\carry[24] ), .Z(SUM[24]) );
  XOR2_X1 U17 ( .A(A[23]), .B(\carry[23] ), .Z(SUM[23]) );
  XOR2_X1 U19 ( .A(A[22]), .B(\carry[22] ), .Z(SUM[22]) );
  XOR2_X1 U21 ( .A(A[21]), .B(\carry[21] ), .Z(SUM[21]) );
  XOR2_X1 U23 ( .A(A[20]), .B(\carry[20] ), .Z(SUM[20]) );
  XOR2_X1 U25 ( .A(A[19]), .B(\carry[19] ), .Z(SUM[19]) );
  XOR2_X1 U27 ( .A(A[18]), .B(\carry[18] ), .Z(SUM[18]) );
  XOR2_X1 U29 ( .A(A[17]), .B(\carry[17] ), .Z(SUM[17]) );
  XOR2_X1 U31 ( .A(A[16]), .B(\carry[16] ), .Z(SUM[16]) );
  XOR2_X1 U33 ( .A(A[15]), .B(\carry[15] ), .Z(SUM[15]) );
  XOR2_X1 U35 ( .A(A[14]), .B(\carry[14] ), .Z(SUM[14]) );
  XOR2_X1 U37 ( .A(A[13]), .B(\carry[13] ), .Z(SUM[13]) );
  XOR2_X1 U39 ( .A(A[12]), .B(\carry[12] ), .Z(SUM[12]) );
  XOR2_X1 U41 ( .A(A[11]), .B(\carry[11] ), .Z(SUM[11]) );
  XOR2_X1 U43 ( .A(A[10]), .B(\carry[10] ), .Z(SUM[10]) );
  XOR2_X1 U45 ( .A(A[9]), .B(\carry[9] ), .Z(SUM[9]) );
  XOR2_X1 U47 ( .A(A[8]), .B(\carry[8] ), .Z(SUM[8]) );
  XOR2_X1 U49 ( .A(A[7]), .B(\carry[7] ), .Z(SUM[7]) );
  XOR2_X1 U51 ( .A(A[6]), .B(\carry[6] ), .Z(SUM[6]) );
  XOR2_X1 U53 ( .A(A[5]), .B(\carry[5] ), .Z(SUM[5]) );
  XOR2_X1 U55 ( .A(A[4]), .B(\carry[4] ), .Z(SUM[4]) );
  XOR2_X1 U57 ( .A(A[3]), .B(\carry[3] ), .Z(SUM[3]) );
  XNOR2_X1 U1 ( .A(A[31]), .B(n1), .ZN(SUM[31]) );
  NAND2_X1 U2 ( .A1(\carry[30] ), .A2(A[30]), .ZN(n1) );
  AND2_X1 U4 ( .A1(\carry[29] ), .A2(A[29]), .ZN(\carry[30] ) );
  AND2_X1 U6 ( .A1(\carry[4] ), .A2(A[4]), .ZN(\carry[5] ) );
  AND2_X1 U8 ( .A1(\carry[5] ), .A2(A[5]), .ZN(\carry[6] ) );
  AND2_X1 U10 ( .A1(\carry[6] ), .A2(A[6]), .ZN(\carry[7] ) );
  AND2_X1 U12 ( .A1(\carry[7] ), .A2(A[7]), .ZN(\carry[8] ) );
  AND2_X1 U14 ( .A1(\carry[8] ), .A2(A[8]), .ZN(\carry[9] ) );
  AND2_X1 U16 ( .A1(\carry[9] ), .A2(A[9]), .ZN(\carry[10] ) );
  AND2_X1 U18 ( .A1(\carry[10] ), .A2(A[10]), .ZN(\carry[11] ) );
  AND2_X1 U20 ( .A1(\carry[11] ), .A2(A[11]), .ZN(\carry[12] ) );
  AND2_X1 U22 ( .A1(\carry[12] ), .A2(A[12]), .ZN(\carry[13] ) );
  AND2_X1 U24 ( .A1(\carry[13] ), .A2(A[13]), .ZN(\carry[14] ) );
  AND2_X1 U26 ( .A1(\carry[14] ), .A2(A[14]), .ZN(\carry[15] ) );
  AND2_X1 U28 ( .A1(\carry[15] ), .A2(A[15]), .ZN(\carry[16] ) );
  AND2_X1 U30 ( .A1(\carry[16] ), .A2(A[16]), .ZN(\carry[17] ) );
  AND2_X1 U32 ( .A1(\carry[17] ), .A2(A[17]), .ZN(\carry[18] ) );
  AND2_X1 U34 ( .A1(\carry[18] ), .A2(A[18]), .ZN(\carry[19] ) );
  AND2_X1 U36 ( .A1(\carry[19] ), .A2(A[19]), .ZN(\carry[20] ) );
  AND2_X1 U38 ( .A1(\carry[20] ), .A2(A[20]), .ZN(\carry[21] ) );
  AND2_X1 U40 ( .A1(\carry[21] ), .A2(A[21]), .ZN(\carry[22] ) );
  AND2_X1 U42 ( .A1(\carry[22] ), .A2(A[22]), .ZN(\carry[23] ) );
  AND2_X1 U44 ( .A1(\carry[23] ), .A2(A[23]), .ZN(\carry[24] ) );
  AND2_X1 U46 ( .A1(\carry[24] ), .A2(A[24]), .ZN(\carry[25] ) );
  AND2_X1 U48 ( .A1(\carry[25] ), .A2(A[25]), .ZN(\carry[26] ) );
  AND2_X1 U50 ( .A1(\carry[26] ), .A2(A[26]), .ZN(\carry[27] ) );
  AND2_X1 U52 ( .A1(\carry[27] ), .A2(A[27]), .ZN(\carry[28] ) );
  AND2_X1 U54 ( .A1(\carry[28] ), .A2(A[28]), .ZN(\carry[29] ) );
  AND2_X1 U56 ( .A1(\carry[3] ), .A2(A[3]), .ZN(\carry[4] ) );
  INV_X1 U58 ( .A(\carry[3] ), .ZN(SUM[2]) );
endmodule


module dlx_cu_FUNC_SIZE11_OP_CODE_SIZE6_CW_SIZE35 ( IR, CLK, RST, RD1_EN, 
        RD2_EN, NPC_LATCH_DEC_EN, REGA_LATCH_EN, REGB_LATCH_EN, 
        REGIMM_LATCH_EN, MUX_SEL_IMM, JUMPFC, MUX_SEL_JAL_ADDR_LW, 
        MUX_SEL_ANPC, MUX_SEL_JAL_IMM, MUX_SEL_BIMM, ALU_OPCODE, 
        MUX_SEL_ALU_32, MUX_SEL_ALU_1, ALU_OUTREG_EN, REGBDELAY_LATCH_EN, 
        DRAM_WE, LMD_LATCH_EN, DRAM_EN, ALU_MA_LATCH_EN, MUX_SEL_WB, RF_WE );
  input [31:0] IR;
  output [1:0] JUMPFC;
  output [1:0] MUX_SEL_JAL_ADDR_LW;
  output [7:0] ALU_OPCODE;
  output [2:0] MUX_SEL_ALU_32;
  output [1:0] MUX_SEL_ALU_1;
  input CLK, RST;
  output RD1_EN, RD2_EN, NPC_LATCH_DEC_EN, REGA_LATCH_EN, REGB_LATCH_EN,
         REGIMM_LATCH_EN, MUX_SEL_IMM, MUX_SEL_ANPC, MUX_SEL_JAL_IMM,
         MUX_SEL_BIMM, ALU_OUTREG_EN, REGBDELAY_LATCH_EN, DRAM_WE,
         LMD_LATCH_EN, DRAM_EN, ALU_MA_LATCH_EN, MUX_SEL_WB, RF_WE;
  wire   IR_31, IR_30, IR_29, IR_28, IR_27, IR_26, cw_15, cw_13, cw_11, cw_10,
         cw_9, cw_8, cw_7, cw_6, cw_5, cw_4, cw_2, cw_0, n30, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n215, n216, n217, n218, n219,
         n220;
  wire   [32:17] cw;
  wire   [23:0] cw1;
  wire   [5:0] cw2;
  wire   [1:0] cw3;
  assign IR_31 = IR[31];
  assign IR_30 = IR[30];
  assign IR_29 = IR[29];
  assign IR_28 = IR[28];
  assign IR_27 = IR[27];
  assign IR_26 = IR[26];
  assign ALU_OPCODE[3] = 1'b0;
  assign MUX_SEL_ALU_32[2] = 1'b0;
  assign RD1_EN = cw[31];

  DFFR_X1 \cw1_reg[32]  ( .D(cw[32]), .CK(CLK), .RN(n215), .Q(NPC_LATCH_DEC_EN) );
  DFFR_X1 \cw1_reg[31]  ( .D(cw[31]), .CK(CLK), .RN(n218), .Q(REGA_LATCH_EN)
         );
  DFFR_X1 \cw1_reg[30]  ( .D(cw[30]), .CK(CLK), .RN(n218), .Q(REGB_LATCH_EN)
         );
  DFFR_X1 \cw1_reg[29]  ( .D(cw[29]), .CK(CLK), .RN(n218), .Q(REGIMM_LATCH_EN)
         );
  DFFR_X1 \cw1_reg[28]  ( .D(cw[28]), .CK(CLK), .RN(n218), .Q(MUX_SEL_IMM) );
  DFFR_X1 \cw1_reg[26]  ( .D(cw[26]), .CK(CLK), .RN(n217), .Q(JUMPFC[0]) );
  DFFR_X1 \cw1_reg[25]  ( .D(cw[25]), .CK(CLK), .RN(n218), .Q(
        MUX_SEL_JAL_ADDR_LW[1]) );
  DFFR_X1 \cw1_reg[24]  ( .D(cw[32]), .CK(CLK), .RN(n215), .Q(
        MUX_SEL_JAL_ADDR_LW[0]) );
  DFFR_X1 \cw1_reg[23]  ( .D(cw[32]), .CK(CLK), .RN(n215), .Q(cw1[23]) );
  DFFR_X1 \cw1_reg[22]  ( .D(cw[31]), .CK(CLK), .RN(n218), .Q(cw1[22]) );
  DFFR_X1 \cw1_reg[21]  ( .D(cw[21]), .CK(CLK), .RN(n218), .Q(cw1[21]) );
  DFFR_X1 \cw1_reg[20]  ( .D(cw[20]), .CK(CLK), .RN(n218), .Q(cw1[20]) );
  DFFR_X1 \cw1_reg[19]  ( .D(cw[19]), .CK(CLK), .RN(n219), .Q(cw1[19]) );
  DFFR_X1 \cw1_reg[18]  ( .D(cw[18]), .CK(CLK), .RN(n219), .Q(cw1[18]) );
  DFFR_X1 \cw1_reg[17]  ( .D(cw[17]), .CK(CLK), .RN(n219), .Q(cw1[17]) );
  DFFR_X1 \cw1_reg[15]  ( .D(cw_15), .CK(CLK), .RN(n216), .Q(cw1[15]) );
  DFFR_X1 \cw1_reg[14]  ( .D(cw_15), .CK(CLK), .RN(n216), .Q(cw1[14]) );
  DFFR_X1 \cw1_reg[13]  ( .D(cw_13), .CK(CLK), .RN(n219), .Q(cw1[13]) );
  DFFR_X1 \cw1_reg[11]  ( .D(cw_11), .CK(CLK), .RN(n219), .Q(cw1[11]) );
  DFFR_X1 \cw1_reg[10]  ( .D(cw_10), .CK(CLK), .RN(n218), .Q(cw1[10]) );
  DFFR_X1 \cw1_reg[9]  ( .D(cw_9), .CK(CLK), .RN(n219), .Q(cw1[9]) );
  DFFR_X1 \cw1_reg[8]  ( .D(cw_8), .CK(CLK), .RN(n219), .Q(cw1[8]) );
  DFFR_X1 \cw1_reg[7]  ( .D(cw_7), .CK(CLK), .RN(n219), .Q(cw1[7]) );
  DFFR_X1 \cw1_reg[6]  ( .D(cw_6), .CK(CLK), .RN(n219), .Q(cw1[6]) );
  DFFR_X1 \cw1_reg[5]  ( .D(cw_5), .CK(CLK), .RN(n217), .Q(cw1[5]) );
  DFFR_X1 \cw1_reg[4]  ( .D(cw_4), .CK(CLK), .RN(n215), .Q(cw1[4]) );
  DFFR_X1 \cw1_reg[3]  ( .D(cw_6), .CK(CLK), .RN(n215), .Q(cw1[3]) );
  DFFR_X1 \cw1_reg[2]  ( .D(cw_2), .CK(CLK), .RN(n215), .Q(cw1[2]) );
  DFFR_X1 \cw1_reg[1]  ( .D(cw_7), .CK(CLK), .RN(n215), .Q(cw1[1]) );
  DFFR_X1 \cw1_reg[0]  ( .D(cw_0), .CK(CLK), .RN(n215), .Q(cw1[0]) );
  DFFR_X1 \cw2_reg[20]  ( .D(cw1[20]), .CK(CLK), .RN(n219), .Q(ALU_OPCODE[7])
         );
  DFFR_X1 \cw2_reg[19]  ( .D(cw1[19]), .CK(CLK), .RN(n219), .Q(ALU_OPCODE[6])
         );
  DFFR_X1 \cw2_reg[18]  ( .D(cw1[18]), .CK(CLK), .RN(n216), .Q(ALU_OPCODE[5])
         );
  DFFR_X1 \cw2_reg[17]  ( .D(cw1[17]), .CK(CLK), .RN(n216), .Q(ALU_OPCODE[4])
         );
  DFFR_X1 \cw2_reg[15]  ( .D(cw1[15]), .CK(CLK), .RN(n216), .Q(ALU_OPCODE[2])
         );
  DFFR_X1 \cw2_reg[14]  ( .D(cw1[14]), .CK(CLK), .RN(n216), .Q(ALU_OPCODE[1])
         );
  DFFR_X1 \cw2_reg[13]  ( .D(cw1[13]), .CK(CLK), .RN(n216), .Q(ALU_OPCODE[0])
         );
  DFFR_X1 \cw2_reg[11]  ( .D(cw1[11]), .CK(CLK), .RN(n216), .Q(
        MUX_SEL_ALU_32[1]) );
  DFFR_X1 \cw2_reg[10]  ( .D(cw1[10]), .CK(CLK), .RN(n219), .Q(
        MUX_SEL_ALU_32[0]) );
  DFFR_X1 \cw2_reg[9]  ( .D(cw1[9]), .CK(CLK), .RN(n216), .Q(MUX_SEL_ALU_1[1])
         );
  DFFR_X1 \cw2_reg[8]  ( .D(cw1[8]), .CK(CLK), .RN(n216), .Q(MUX_SEL_ALU_1[0])
         );
  DFFR_X1 \cw2_reg[7]  ( .D(cw1[7]), .CK(CLK), .RN(n216), .Q(ALU_OUTREG_EN) );
  DFFR_X1 \cw2_reg[6]  ( .D(cw1[6]), .CK(CLK), .RN(n216), .Q(
        REGBDELAY_LATCH_EN) );
  DFFR_X1 \cw2_reg[5]  ( .D(cw1[5]), .CK(CLK), .RN(n218), .Q(cw2[5]) );
  DFFR_X1 \cw2_reg[4]  ( .D(cw1[4]), .CK(CLK), .RN(n217), .Q(cw2[4]) );
  DFFR_X1 \cw2_reg[3]  ( .D(cw1[3]), .CK(CLK), .RN(n217), .Q(cw2[3]) );
  DFFR_X1 \cw2_reg[2]  ( .D(cw1[2]), .CK(CLK), .RN(n217), .Q(cw2[2]) );
  DFFR_X1 \cw2_reg[1]  ( .D(cw1[1]), .CK(CLK), .RN(n217), .Q(cw2[1]) );
  DFFR_X1 \cw2_reg[0]  ( .D(cw1[0]), .CK(CLK), .RN(n217), .Q(cw2[0]) );
  DFFR_X1 \cw3_reg[5]  ( .D(cw2[5]), .CK(CLK), .RN(n218), .Q(DRAM_WE) );
  DFFR_X1 \cw3_reg[4]  ( .D(cw2[4]), .CK(CLK), .RN(n217), .Q(LMD_LATCH_EN) );
  DFFR_X1 \cw3_reg[3]  ( .D(cw2[3]), .CK(CLK), .RN(n217), .Q(DRAM_EN) );
  DFFR_X1 \cw3_reg[2]  ( .D(cw2[2]), .CK(CLK), .RN(n215), .Q(ALU_MA_LATCH_EN)
         );
  DFFR_X1 \cw3_reg[1]  ( .D(cw2[1]), .CK(CLK), .RN(n217), .Q(cw3[1]) );
  DFFR_X1 \cw4_reg[1]  ( .D(cw3[1]), .CK(CLK), .RN(n217), .Q(MUX_SEL_WB) );
  DFFR_X1 \cw3_reg[0]  ( .D(cw2[0]), .CK(CLK), .RN(n215), .Q(cw3[0]) );
  DFFR_X1 \cw4_reg[0]  ( .D(cw3[0]), .CK(CLK), .RN(n218), .Q(RF_WE) );
  DFFR_X1 \cw1_reg[27]  ( .D(n30), .CK(CLK), .RN(n217), .Q(JUMPFC[1]) );
  DFFR_X1 \cw2_reg[23]  ( .D(cw1[23]), .CK(CLK), .RN(n220), .Q(MUX_SEL_ANPC)
         );
  DFFR_X1 \cw2_reg[22]  ( .D(cw1[22]), .CK(CLK), .RN(n215), .Q(MUX_SEL_JAL_IMM) );
  DFFR_X1 \cw2_reg[21]  ( .D(cw1[21]), .CK(CLK), .RN(n215), .Q(MUX_SEL_BIMM)
         );
  OAI33_X1 U85 ( .A1(n88), .A2(n89), .A3(n90), .B1(n91), .B2(n92), .B3(n93), 
        .ZN(cw_8) );
  NAND3_X1 U86 ( .A1(IR_27), .A2(IR_28), .A3(n110), .ZN(n109) );
  OAI33_X1 U87 ( .A1(n91), .A2(IR_30), .A3(n92), .B1(n112), .B2(n113), .B3(
        n114), .ZN(n111) );
  NAND3_X1 U88 ( .A1(n116), .A2(n117), .A3(n118), .ZN(cw_2) );
  NAND3_X1 U89 ( .A1(n131), .A2(n102), .A3(n128), .ZN(cw[18]) );
  NAND3_X1 U90 ( .A1(n136), .A2(n137), .A3(n107), .ZN(cw[17]) );
  OAI33_X1 U91 ( .A1(n93), .A2(IR_26), .A3(n92), .B1(n139), .B2(IR[1]), .B3(
        n140), .ZN(cw_9) );
  NAND3_X1 U92 ( .A1(IR_30), .A2(n141), .A3(IR_26), .ZN(n100) );
  NAND3_X1 U93 ( .A1(IR_27), .A2(n134), .A3(n110), .ZN(n136) );
  NAND3_X1 U94 ( .A1(n119), .A2(n142), .A3(IR_31), .ZN(n115) );
  NAND3_X1 U95 ( .A1(n134), .A2(n93), .A3(IR_27), .ZN(n124) );
  NAND3_X1 U96 ( .A1(n91), .A2(n134), .A3(n146), .ZN(n89) );
  NAND3_X1 U97 ( .A1(n143), .A2(n149), .A3(IR[2]), .ZN(n147) );
  INV_X1 U5 ( .A(n121), .ZN(cw[30]) );
  NOR2_X1 U6 ( .A1(cw[21]), .A2(cw_6), .ZN(n121) );
  INV_X1 U7 ( .A(n89), .ZN(n104) );
  NAND2_X1 U8 ( .A1(n135), .A2(n104), .ZN(n112) );
  NAND2_X1 U9 ( .A1(n118), .A2(n121), .ZN(cw[31]) );
  INV_X1 U10 ( .A(cw_2), .ZN(n94) );
  INV_X1 U11 ( .A(n95), .ZN(cw_6) );
  NAND2_X1 U12 ( .A1(n94), .A2(n95), .ZN(cw_7) );
  NAND2_X1 U13 ( .A1(n118), .A2(n95), .ZN(cw[29]) );
  OR2_X1 U14 ( .A1(n30), .A2(cw[31]), .ZN(cw[28]) );
  INV_X1 U15 ( .A(n117), .ZN(cw[32]) );
  NOR3_X1 U16 ( .A1(n134), .A2(n123), .A3(n93), .ZN(n133) );
  NOR2_X1 U17 ( .A1(cw_4), .A2(cw_5), .ZN(n95) );
  OAI21_X1 U18 ( .B1(n147), .B2(n148), .A(n88), .ZN(n105) );
  NAND2_X1 U19 ( .A1(n114), .A2(n113), .ZN(n148) );
  AOI21_X1 U20 ( .B1(n113), .B2(n108), .A(n106), .ZN(n128) );
  NOR2_X1 U21 ( .A1(n124), .A2(n91), .ZN(n119) );
  OR4_X1 U22 ( .A1(n114), .A2(n149), .A3(n113), .A4(n150), .ZN(n88) );
  INV_X1 U23 ( .A(cw_9), .ZN(n101) );
  AND3_X1 U24 ( .A1(n125), .A2(n102), .A3(n126), .ZN(n118) );
  AND3_X1 U25 ( .A1(n100), .A2(n127), .A3(n92), .ZN(n126) );
  INV_X1 U26 ( .A(n110), .ZN(n127) );
  NAND2_X1 U27 ( .A1(n133), .A2(IR_27), .ZN(n102) );
  OAI21_X1 U28 ( .B1(n96), .B2(n97), .A(n98), .ZN(cw_15) );
  INV_X1 U29 ( .A(n143), .ZN(n150) );
  NAND4_X1 U30 ( .A1(n100), .A2(n101), .A3(n102), .A4(n103), .ZN(cw_11) );
  AOI21_X1 U31 ( .B1(n104), .B2(n105), .A(n106), .ZN(n103) );
  INV_X1 U32 ( .A(n147), .ZN(n135) );
  INV_X1 U33 ( .A(n120), .ZN(n123) );
  INV_X1 U34 ( .A(n115), .ZN(cw_4) );
  NAND4_X1 U35 ( .A1(n107), .A2(n98), .A3(n92), .A4(n96), .ZN(cw_10) );
  INV_X1 U36 ( .A(n106), .ZN(n125) );
  NAND2_X1 U37 ( .A1(n118), .A2(n115), .ZN(cw[25]) );
  NAND2_X1 U38 ( .A1(n115), .A2(n94), .ZN(cw_0) );
  INV_X1 U39 ( .A(n138), .ZN(n107) );
  OAI211_X1 U40 ( .C1(n89), .C2(n88), .A(n100), .B(n101), .ZN(n138) );
  INV_X1 U41 ( .A(n116), .ZN(cw[21]) );
  OAI21_X1 U42 ( .B1(n129), .B2(n130), .A(n125), .ZN(cw[19]) );
  NAND2_X1 U43 ( .A1(n97), .A2(n113), .ZN(n130) );
  INV_X1 U44 ( .A(n108), .ZN(n129) );
  OAI22_X1 U45 ( .A1(n91), .A2(n122), .B1(n123), .B2(n124), .ZN(cw[26]) );
  NAND2_X1 U46 ( .A1(n119), .A2(n120), .ZN(n117) );
  INV_X1 U47 ( .A(n122), .ZN(n30) );
  NAND2_X1 U48 ( .A1(IR[3]), .A2(IR[2]), .ZN(n139) );
  NOR4_X1 U49 ( .A1(IR[6]), .A2(IR[4]), .A3(IR[10]), .A4(n153), .ZN(n143) );
  OR3_X1 U50 ( .A1(IR[9]), .A2(IR[8]), .A3(IR[7]), .ZN(n153) );
  NOR4_X1 U51 ( .A1(n142), .A2(IR_26), .A3(IR_30), .A4(IR_31), .ZN(n110) );
  INV_X1 U52 ( .A(IR[2]), .ZN(n90) );
  NOR3_X1 U53 ( .A1(IR_26), .A2(IR_27), .A3(n132), .ZN(n106) );
  INV_X1 U54 ( .A(n133), .ZN(n132) );
  NOR3_X1 U55 ( .A1(IR_27), .A2(IR_30), .A3(n123), .ZN(n146) );
  NOR3_X1 U56 ( .A1(IR_27), .A2(IR_31), .A3(n142), .ZN(n141) );
  NOR2_X1 U57 ( .A1(n112), .A2(IR[0]), .ZN(n108) );
  OAI221_X1 U58 ( .B1(IR[1]), .B2(n96), .C1(IR_30), .C2(n92), .A(n99), .ZN(
        cw_13) );
  INV_X1 U59 ( .A(IR[1]), .ZN(n97) );
  INV_X1 U60 ( .A(IR[5]), .ZN(n113) );
  NOR2_X1 U61 ( .A1(IR_29), .A2(IR_31), .ZN(n120) );
  NAND4_X1 U62 ( .A1(IR[5]), .A2(n143), .A3(n104), .A4(n144), .ZN(n140) );
  NAND2_X1 U63 ( .A1(n141), .A2(IR_28), .ZN(n92) );
  OAI21_X1 U64 ( .B1(n145), .B2(n105), .A(n104), .ZN(n116) );
  NOR4_X1 U65 ( .A1(n151), .A2(n152), .A3(n150), .A4(n113), .ZN(n145) );
  AOI21_X1 U66 ( .B1(IR[2]), .B2(n97), .A(n149), .ZN(n152) );
  AOI21_X1 U67 ( .B1(n135), .B2(n97), .A(n144), .ZN(n151) );
  NAND2_X1 U68 ( .A1(n108), .A2(IR[5]), .ZN(n96) );
  INV_X1 U69 ( .A(IR_26), .ZN(n91) );
  NAND2_X1 U70 ( .A1(IR_28), .A2(n146), .ZN(n122) );
  INV_X1 U71 ( .A(n111), .ZN(n99) );
  INV_X1 U72 ( .A(IR_30), .ZN(n93) );
  OAI21_X1 U73 ( .B1(IR_26), .B2(n102), .A(n128), .ZN(cw[20]) );
  NAND2_X1 U74 ( .A1(IR[0]), .A2(n97), .ZN(n114) );
  INV_X1 U75 ( .A(IR_28), .ZN(n134) );
  INV_X1 U76 ( .A(IR_29), .ZN(n142) );
  AND2_X1 U77 ( .A1(n99), .A2(n109), .ZN(n98) );
  AND3_X1 U78 ( .A1(n119), .A2(IR_29), .A3(IR_31), .ZN(cw_5) );
  INV_X1 U79 ( .A(IR[0]), .ZN(n144) );
  OR3_X1 U80 ( .A1(n112), .A2(IR[5]), .A3(n97), .ZN(n131) );
  INV_X1 U81 ( .A(IR[3]), .ZN(n149) );
  OR4_X1 U82 ( .A1(n97), .A2(n140), .A3(IR[2]), .A4(IR[3]), .ZN(n137) );
  NAND2_X1 U83 ( .A1(n122), .A2(n121), .ZN(RD2_EN) );
  CLKBUF_X1 U84 ( .A(n220), .Z(n215) );
  CLKBUF_X1 U98 ( .A(n220), .Z(n216) );
  CLKBUF_X1 U99 ( .A(n220), .Z(n217) );
  CLKBUF_X1 U100 ( .A(n220), .Z(n218) );
  CLKBUF_X1 U101 ( .A(n220), .Z(n219) );
  INV_X1 U102 ( .A(RST), .ZN(n220) );
endmodule


module datapath ( CLK, RST, SOURCE1, SOURCE2, DESTINATION, IMMEDIATE, NPC, 
        RD1_EN, RD2_EN, REGA_LATCH_EN, REGB_LATCH_EN, REGIMM_LATCH_EN, 
        MUX_SEL_IMM, MUX_SEL_JAL_ADDR_LW, NPC_LATCH_DEC_EN, JUMPFC, 
        NPC_DATAPATH_OUT, REG_DELAY1, REG_DELAY2, REG_DELAY3, REG_DELAY4, 
        EN_IN, ALU_OPCODE, MUX_SEL_JAL_IMM, MUX_SEL_BIMM, MUX_SEL_ANPC, 
        MUX_SEL_ALU_32, MUX_SEL_ALU_1, ALU_OUTREG_EN, REGBDELAY_LATCH_EN, 
        DRAM_WE, LMD_LATCH_EN, ALU_MA_LATCH_EN, DRAM_EN, MUX_SEL_WB, RF_WE );
  input [4:0] SOURCE1;
  input [4:0] SOURCE2;
  input [5:0] DESTINATION;
  input [25:0] IMMEDIATE;
  input [31:0] NPC;
  input [1:0] MUX_SEL_JAL_ADDR_LW;
  input [1:0] JUMPFC;
  output [31:0] NPC_DATAPATH_OUT;
  output [5:0] REG_DELAY1;
  output [5:0] REG_DELAY2;
  output [5:0] REG_DELAY3;
  output [5:0] REG_DELAY4;
  input [7:0] ALU_OPCODE;
  input [2:0] MUX_SEL_ALU_32;
  input [1:0] MUX_SEL_ALU_1;
  input CLK, RST, RD1_EN, RD2_EN, REGA_LATCH_EN, REGB_LATCH_EN,
         REGIMM_LATCH_EN, MUX_SEL_IMM, NPC_LATCH_DEC_EN, EN_IN,
         MUX_SEL_JAL_IMM, MUX_SEL_BIMM, MUX_SEL_ANPC, ALU_OUTREG_EN,
         REGBDELAY_LATCH_EN, DRAM_WE, LMD_LATCH_EN, ALU_MA_LATCH_EN, DRAM_EN,
         MUX_SEL_WB, RF_WE;
  wire   sig_flush;
  wire   [31:0] sig_rf_datain;
  wire   [31:0] sig_rega;
  wire   [31:0] sig_regb_decode;
  wire   [31:0] sig_imm;
  wire   [31:0] sig_npc_ex_in;
  wire   [31:0] sig_regalu;
  wire   [31:0] sig_regb_ex;
  wire   [31:0] sig_alu_ma;
  wire   [31:0] sig_lmd;

  decode_stage decode_map ( .RST(RST), .CLK(CLK), .SOURCE1(SOURCE1), .SOURCE2(
        SOURCE2), .DESTINATION(DESTINATION), .IMMEDIATE(IMMEDIATE), .NPC(NPC), 
        .RD1_EN(RD1_EN), .RD2_EN(RD2_EN), .WR_EN_WB(RF_WE), .RF_DATAIN(
        sig_rf_datain), .REGA_LATCH_EN(REGA_LATCH_EN), .REGB_LATCH_EN(
        REGB_LATCH_EN), .REGIMM_LATCH_EN(REGIMM_LATCH_EN), .NPC_LATCH_DEC_EN(
        NPC_LATCH_DEC_EN), .MUX_SEL_IMM(MUX_SEL_IMM), .JUMPFC(JUMPFC), 
        .MUX_SEL_JAL_ADDR_LW(MUX_SEL_JAL_ADDR_LW), .REGA_OUT(sig_rega), 
        .REGB_OUT(sig_regb_decode), .REGIMM_OUT(sig_imm), .NPC_EXECUTE_IN(
        sig_npc_ex_in), .NPC_DECODE_OUT(NPC_DATAPATH_OUT), .FLUSH(sig_flush), 
        .REG_DELAY1(REG_DELAY1), .REG_DELAY2(REG_DELAY2), .REG_DELAY3(
        REG_DELAY3), .REG_DELAY4(REG_DELAY4), .EN_IN(EN_IN) );
  execute_stage execute_map ( .CLK(CLK), .RST(RST), .NPC_EXECUTE_IN(
        sig_npc_ex_in), .REGA_OUT(sig_rega), .REGB_OUT(sig_regb_decode), 
        .REGIMM_OUT(sig_imm), .ALU_OPCODE(ALU_OPCODE), .MUX_SEL_ANPC(
        MUX_SEL_ANPC), .MUX_SEL_BIMM(MUX_SEL_BIMM), .MUX_SEL_JAL_IMM(
        MUX_SEL_JAL_IMM), .MUX_SEL_ALU_32(MUX_SEL_ALU_32), .MUX_SEL_ALU_1(
        MUX_SEL_ALU_1), .ALU_OUTREG_EN(ALU_OUTREG_EN), .REGBDELAY_LATCH_EN(
        REGBDELAY_LATCH_EN), .REGALU_OUT(sig_regalu), .REGB_EX_OUT(sig_regb_ex) );
  mem_access_stage mem_access_map ( .ALU_OUT(sig_regalu), .REGB_EX_OUT(
        sig_regb_ex), .DRAM_WE(DRAM_WE), .LMD_LATCH_EN(LMD_LATCH_EN), 
        .DRAM_EN(DRAM_EN), .RST(RST), .CLK(CLK), .ALU_MA_LATCH_EN(
        ALU_MA_LATCH_EN), .FLUSH(sig_flush), .ALU_MA_OUT(sig_alu_ma), 
        .LMD_OUT(sig_lmd) );
  write_back_stage write_back_map ( .LMD_OUT(sig_lmd), .ALU_MA_OUT(sig_alu_ma), 
        .MUX_SEL_WB(MUX_SEL_WB), .RF_DATA_IN(sig_rf_datain) );
endmodule


module dependency_manager ( RST, IR, IR_OUT, DIRTY_BIT, EN_OUT, REG_DELAY1, 
        REG_DELAY2, REG_DELAY3, REG_DELAY4 );
  input [31:0] IR;
  output [31:0] IR_OUT;
  input [5:0] REG_DELAY1;
  input [5:0] REG_DELAY2;
  input [5:0] REG_DELAY3;
  input [5:0] REG_DELAY4;
  input RST;
  output DIRTY_BIT, EN_OUT;
  wire   N496, n128, n11, n12, n13, n14, n15, n16, n17, n18, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n123, n124, n126, n127;

  DLL_X1 DIRTY_BIT_reg ( .D(N496), .GN(RST), .Q(DIRTY_BIT) );
  XOR2_X1 U82 ( .A(REG_DELAY3[0]), .B(IR[16]), .Z(n35) );
  XOR2_X1 U83 ( .A(REG_DELAY3[4]), .B(IR[20]), .Z(n34) );
  XOR2_X1 U84 ( .A(REG_DELAY3[1]), .B(IR[17]), .Z(n33) );
  XOR2_X1 U88 ( .A(REG_DELAY2[1]), .B(IR[17]), .Z(n44) );
  XOR2_X1 U89 ( .A(REG_DELAY2[4]), .B(IR[20]), .Z(n43) );
  XOR2_X1 U90 ( .A(REG_DELAY2[3]), .B(n21), .Z(n41) );
  XOR2_X1 U91 ( .A(REG_DELAY2[2]), .B(n22), .Z(n40) );
  XOR2_X1 U92 ( .A(REG_DELAY2[0]), .B(n24), .Z(n39) );
  XOR2_X1 U93 ( .A(REG_DELAY4[1]), .B(IR[17]), .Z(n50) );
  XOR2_X1 U94 ( .A(REG_DELAY4[4]), .B(IR[20]), .Z(n49) );
  XOR2_X1 U95 ( .A(REG_DELAY4[3]), .B(n21), .Z(n47) );
  XOR2_X1 U96 ( .A(REG_DELAY4[2]), .B(n22), .Z(n46) );
  XOR2_X1 U97 ( .A(REG_DELAY4[0]), .B(n24), .Z(n45) );
  XOR2_X1 U98 ( .A(REG_DELAY1[2]), .B(IR[18]), .Z(n56) );
  XOR2_X1 U99 ( .A(REG_DELAY1[3]), .B(IR[19]), .Z(n55) );
  XOR2_X1 U100 ( .A(REG_DELAY1[1]), .B(n23), .Z(n53) );
  XOR2_X1 U101 ( .A(REG_DELAY1[0]), .B(n24), .Z(n52) );
  XOR2_X1 U102 ( .A(REG_DELAY1[4]), .B(n20), .Z(n51) );
  XOR2_X1 U103 ( .A(REG_DELAY2[1]), .B(IR[22]), .Z(n66) );
  XOR2_X1 U104 ( .A(REG_DELAY2[4]), .B(IR[25]), .Z(n65) );
  XOR2_X1 U105 ( .A(REG_DELAY1[1]), .B(IR[22]), .Z(n72) );
  XOR2_X1 U106 ( .A(REG_DELAY1[4]), .B(IR[25]), .Z(n71) );
  XOR2_X1 U107 ( .A(REG_DELAY4[1]), .B(IR[22]), .Z(n78) );
  XOR2_X1 U108 ( .A(REG_DELAY4[4]), .B(IR[25]), .Z(n77) );
  XOR2_X1 U109 ( .A(REG_DELAY3[1]), .B(IR[22]), .Z(n84) );
  XOR2_X1 U110 ( .A(REG_DELAY3[4]), .B(IR[25]), .Z(n83) );
  INV_X1 U3 ( .A(n127), .ZN(n126) );
  INV_X1 U4 ( .A(n15), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n127), .A2(n16), .ZN(IR_OUT[27]) );
  NAND4_X1 U6 ( .A1(n57), .A2(n58), .A3(n59), .A4(n60), .ZN(n15) );
  NAND4_X1 U7 ( .A1(n79), .A2(n80), .A3(n81), .A4(n82), .ZN(n57) );
  NAND4_X1 U8 ( .A1(n73), .A2(n74), .A3(n75), .A4(n76), .ZN(n58) );
  NAND4_X1 U9 ( .A1(n67), .A2(n68), .A3(n69), .A4(n70), .ZN(n59) );
  INV_X1 U10 ( .A(n11), .ZN(n17) );
  AND4_X1 U11 ( .A1(n27), .A2(n28), .A3(n29), .A4(n30), .ZN(n18) );
  NAND4_X1 U12 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(n27) );
  NAND4_X1 U13 ( .A1(n45), .A2(n46), .A3(n47), .A4(n48), .ZN(n28) );
  NAND4_X1 U14 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(n29) );
  NOR2_X1 U15 ( .A1(n127), .A2(n21), .ZN(IR_OUT[19]) );
  NOR2_X1 U16 ( .A1(n127), .A2(n24), .ZN(IR_OUT[16]) );
  NOR2_X1 U17 ( .A1(n127), .A2(n20), .ZN(IR_OUT[20]) );
  NOR2_X1 U18 ( .A1(n127), .A2(n23), .ZN(IR_OUT[17]) );
  NOR2_X1 U19 ( .A1(n127), .A2(n22), .ZN(IR_OUT[18]) );
  NOR4_X1 U20 ( .A1(IR[28]), .A2(IR[29]), .A3(IR[30]), .A4(IR[31]), .ZN(n11)
         );
  NOR3_X1 U21 ( .A1(n43), .A2(REG_DELAY2[5]), .A3(n44), .ZN(n42) );
  NOR3_X1 U22 ( .A1(n49), .A2(REG_DELAY4[5]), .A3(n50), .ZN(n48) );
  NOR3_X1 U23 ( .A1(n55), .A2(REG_DELAY1[5]), .A3(n56), .ZN(n54) );
  NOR3_X1 U24 ( .A1(n71), .A2(REG_DELAY1[5]), .A3(n72), .ZN(n70) );
  NOR3_X1 U25 ( .A1(n77), .A2(REG_DELAY4[5]), .A3(n78), .ZN(n76) );
  NOR3_X1 U26 ( .A1(n83), .A2(REG_DELAY3[5]), .A3(n84), .ZN(n82) );
  NOR3_X1 U27 ( .A1(n65), .A2(REG_DELAY2[5]), .A3(n66), .ZN(n64) );
  AND2_X1 U28 ( .A1(n126), .A2(IR[25]), .ZN(IR_OUT[25]) );
  AND2_X1 U29 ( .A1(n126), .A2(IR[21]), .ZN(IR_OUT[21]) );
  AND2_X1 U30 ( .A1(n126), .A2(IR[24]), .ZN(IR_OUT[24]) );
  AND2_X1 U31 ( .A1(n126), .A2(IR[30]), .ZN(IR_OUT[30]) );
  AND2_X1 U32 ( .A1(n126), .A2(IR[26]), .ZN(IR_OUT[26]) );
  OR3_X1 U33 ( .A1(n123), .A2(REG_DELAY3[5]), .A3(n124), .ZN(n32) );
  XNOR2_X1 U34 ( .A(REG_DELAY3[3]), .B(n21), .ZN(n123) );
  XNOR2_X1 U35 ( .A(REG_DELAY3[2]), .B(n22), .ZN(n124) );
  AND2_X1 U36 ( .A1(n126), .A2(IR[31]), .ZN(IR_OUT[31]) );
  AND2_X1 U37 ( .A1(IR[2]), .A2(n126), .ZN(IR_OUT[2]) );
  AND2_X1 U38 ( .A1(IR[5]), .A2(n126), .ZN(IR_OUT[5]) );
  XNOR2_X1 U39 ( .A(REG_DELAY1[3]), .B(IR[24]), .ZN(n69) );
  XNOR2_X1 U40 ( .A(REG_DELAY4[3]), .B(IR[24]), .ZN(n75) );
  XNOR2_X1 U41 ( .A(REG_DELAY3[3]), .B(IR[24]), .ZN(n81) );
  XNOR2_X1 U42 ( .A(REG_DELAY1[2]), .B(IR[23]), .ZN(n68) );
  XNOR2_X1 U43 ( .A(REG_DELAY4[2]), .B(IR[23]), .ZN(n74) );
  XNOR2_X1 U44 ( .A(REG_DELAY3[2]), .B(IR[23]), .ZN(n80) );
  AND2_X1 U45 ( .A1(n126), .A2(IR[28]), .ZN(IR_OUT[28]) );
  AND2_X1 U46 ( .A1(IR[0]), .A2(EN_OUT), .ZN(IR_OUT[0]) );
  NOR2_X1 U47 ( .A1(n31), .A2(n15), .ZN(n30) );
  NOR4_X1 U48 ( .A1(n32), .A2(n33), .A3(n34), .A4(n35), .ZN(n31) );
  NAND4_X1 U49 ( .A1(n61), .A2(n62), .A3(n63), .A4(n64), .ZN(n60) );
  XNOR2_X1 U50 ( .A(REG_DELAY2[0]), .B(IR[21]), .ZN(n61) );
  XNOR2_X1 U51 ( .A(REG_DELAY2[2]), .B(IR[23]), .ZN(n62) );
  XNOR2_X1 U52 ( .A(REG_DELAY2[3]), .B(IR[24]), .ZN(n63) );
  AND2_X1 U53 ( .A1(n126), .A2(IR[23]), .ZN(IR_OUT[23]) );
  XNOR2_X1 U54 ( .A(REG_DELAY1[0]), .B(IR[21]), .ZN(n67) );
  XNOR2_X1 U55 ( .A(REG_DELAY4[0]), .B(IR[21]), .ZN(n73) );
  XNOR2_X1 U56 ( .A(REG_DELAY3[0]), .B(IR[21]), .ZN(n79) );
  INV_X1 U57 ( .A(IR[19]), .ZN(n21) );
  INV_X1 U58 ( .A(IR[18]), .ZN(n22) );
  INV_X1 U59 ( .A(IR[16]), .ZN(n24) );
  OAI211_X1 U60 ( .C1(n17), .C2(n16), .A(n25), .B(n26), .ZN(n128) );
  OAI21_X1 U61 ( .B1(IR[26]), .B2(n17), .A(n12), .ZN(n25) );
  NOR2_X1 U62 ( .A1(RST), .A2(n18), .ZN(n26) );
  AND2_X1 U63 ( .A1(IR[1]), .A2(n126), .ZN(IR_OUT[1]) );
  AND2_X1 U64 ( .A1(n126), .A2(IR[22]), .ZN(IR_OUT[22]) );
  AND2_X1 U65 ( .A1(IR[3]), .A2(n126), .ZN(IR_OUT[3]) );
  AND2_X1 U66 ( .A1(n126), .A2(IR[29]), .ZN(IR_OUT[29]) );
  INV_X1 U67 ( .A(IR[27]), .ZN(n16) );
  AND2_X1 U68 ( .A1(IR[7]), .A2(EN_OUT), .ZN(IR_OUT[7]) );
  AND2_X1 U69 ( .A1(IR[8]), .A2(EN_OUT), .ZN(IR_OUT[8]) );
  INV_X1 U70 ( .A(IR[17]), .ZN(n23) );
  INV_X1 U71 ( .A(IR[20]), .ZN(n20) );
  AND2_X1 U72 ( .A1(IR[10]), .A2(n126), .ZN(IR_OUT[10]) );
  AND2_X1 U73 ( .A1(IR[4]), .A2(n126), .ZN(IR_OUT[4]) );
  AND2_X1 U74 ( .A1(IR[6]), .A2(n126), .ZN(IR_OUT[6]) );
  AND2_X1 U75 ( .A1(IR[9]), .A2(n126), .ZN(IR_OUT[9]) );
  OAI21_X1 U76 ( .B1(n11), .B2(n12), .A(n13), .ZN(N496) );
  OAI21_X1 U77 ( .B1(n14), .B2(n15), .A(n16), .ZN(n13) );
  NOR3_X1 U78 ( .A1(n17), .A2(IR[26]), .A3(n18), .ZN(n14) );
  AND2_X1 U79 ( .A1(IR[11]), .A2(n126), .ZN(IR_OUT[11]) );
  AND2_X1 U80 ( .A1(IR[12]), .A2(n126), .ZN(IR_OUT[12]) );
  AND2_X1 U81 ( .A1(IR[13]), .A2(n126), .ZN(IR_OUT[13]) );
  AND2_X1 U85 ( .A1(IR[14]), .A2(n126), .ZN(IR_OUT[14]) );
  AND2_X1 U86 ( .A1(IR[15]), .A2(n126), .ZN(IR_OUT[15]) );
  INV_X1 U87 ( .A(n127), .ZN(EN_OUT) );
  INV_X1 U111 ( .A(n128), .ZN(n127) );
endmodule


module Add4_N32 ( A, Y );
  input [31:0] A;
  output [31:0] Y;


  Add4_N32_DW01_add_0 add_17 ( .A(A), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b0, 1'b0}), .CI(1'b0), .SUM(Y) );
endmodule


module reg_generic_N32 ( D, CLK, RST, EN, Q );
  input [31:0] D;
  output [31:0] Q;
  input CLK, RST, EN;
  wire   n6, n7;
  assign n6 = RST;
  assign n7 = EN;

  FD_s_0 UFD_0 ( .D(D[0]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[0]) );
  FD_s_31 UFD_1 ( .D(D[1]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[1]) );
  FD_s_30 UFD_2 ( .D(D[2]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[2]) );
  FD_s_29 UFD_3 ( .D(D[3]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[3]) );
  FD_s_28 UFD_4 ( .D(D[4]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[4]) );
  FD_s_27 UFD_5 ( .D(D[5]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[5]) );
  FD_s_26 UFD_6 ( .D(D[6]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[6]) );
  FD_s_25 UFD_7 ( .D(D[7]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[7]) );
  FD_s_24 UFD_8 ( .D(D[8]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[8]) );
  FD_s_23 UFD_9 ( .D(D[9]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[9]) );
  FD_s_22 UFD_10 ( .D(D[10]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[10]) );
  FD_s_21 UFD_11 ( .D(D[11]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[11]) );
  FD_s_20 UFD_12 ( .D(D[12]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[12]) );
  FD_s_19 UFD_13 ( .D(D[13]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[13]) );
  FD_s_18 UFD_14 ( .D(D[14]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[14]) );
  FD_s_17 UFD_15 ( .D(D[15]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[15]) );
  FD_s_16 UFD_16 ( .D(D[16]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[16]) );
  FD_s_15 UFD_17 ( .D(D[17]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[17]) );
  FD_s_14 UFD_18 ( .D(D[18]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[18]) );
  FD_s_13 UFD_19 ( .D(D[19]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[19]) );
  FD_s_12 UFD_20 ( .D(D[20]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[20]) );
  FD_s_11 UFD_21 ( .D(D[21]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[21]) );
  FD_s_10 UFD_22 ( .D(D[22]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[22]) );
  FD_s_9 UFD_23 ( .D(D[23]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[23]) );
  FD_s_8 UFD_24 ( .D(D[24]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[24]) );
  FD_s_7 UFD_25 ( .D(D[25]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[25]) );
  FD_s_6 UFD_26 ( .D(D[26]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[26]) );
  FD_s_5 UFD_27 ( .D(D[27]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[27]) );
  FD_s_4 UFD_28 ( .D(D[28]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[28]) );
  FD_s_3 UFD_29 ( .D(D[29]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[29]) );
  FD_s_2 UFD_30 ( .D(D[30]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[30]) );
  FD_s_1 UFD_31 ( .D(D[31]), .CLK(CLK), .RST(n6), .EN(n7), .Q(Q[31]) );
endmodule


module top_entity ( CLK, RST, PC, IR );
  output [31:0] PC;
  input [31:0] IR;
  input CLK, RST;
  wire   sig_en_dependecy, \sig_destination[5] , sig_rd1_en, sig_rd2_en,
         sig_rega_latch_en, sig_regb_latch_en, sig_regimm_latch_en,
         sig_mux_sel_imm, sig_npc_latch_dec_en, sig_mux_sel_jal_imm,
         sig_mux_sel_bimm, sig_sel_anpc, sig_alu_outreg_en,
         sig_regbdelay_latch_en, sig_dram_we, sig_lmd_latch_en,
         sig_alu_ma_latch_en, sig_dram_en, sig_mux_sel_wb, sig_rf_we;
  wire   [31:0] sig_npc_datapath;
  wire   [31:0] sig_npc;
  wire   [31:0] sig_ir_dependency;
  wire   [5:0] sig_reg_delay1;
  wire   [5:0] sig_reg_delay2;
  wire   [5:0] sig_reg_delay3;
  wire   [5:0] sig_reg_delay4;
  wire   [1:0] sig_mux_sel_jal_addr;
  wire   [1:0] sig_jumpfc;
  wire   [7:0] sig_alu_opcode;
  wire   [2:0] sig_mux_sel_alu_32;
  wire   [1:0] sig_mux_sel_alu_1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  reg_generic_N32 reg_pc ( .D(sig_npc_datapath), .CLK(CLK), .RST(RST), .EN(
        sig_en_dependecy), .Q(PC) );
  Add4_N32 add4_0 ( .A(PC), .Y(sig_npc) );
  dependency_manager dep_man ( .RST(RST), .IR(IR), .IR_OUT(sig_ir_dependency), 
        .DIRTY_BIT(\sig_destination[5] ), .EN_OUT(sig_en_dependecy), 
        .REG_DELAY1(sig_reg_delay1), .REG_DELAY2(sig_reg_delay2), .REG_DELAY3(
        sig_reg_delay3), .REG_DELAY4(sig_reg_delay4) );
  datapath datapath_0 ( .CLK(CLK), .RST(RST), .SOURCE1(
        sig_ir_dependency[25:21]), .SOURCE2(sig_ir_dependency[20:16]), 
        .DESTINATION({\sig_destination[5] , sig_ir_dependency[15:11]}), 
        .IMMEDIATE(sig_ir_dependency[25:0]), .NPC(sig_npc), .RD1_EN(sig_rd1_en), .RD2_EN(sig_rd2_en), .REGA_LATCH_EN(sig_rega_latch_en), .REGB_LATCH_EN(
        sig_regb_latch_en), .REGIMM_LATCH_EN(sig_regimm_latch_en), 
        .MUX_SEL_IMM(sig_mux_sel_imm), .MUX_SEL_JAL_ADDR_LW(
        sig_mux_sel_jal_addr), .NPC_LATCH_DEC_EN(sig_npc_latch_dec_en), 
        .JUMPFC(sig_jumpfc), .NPC_DATAPATH_OUT(sig_npc_datapath), .REG_DELAY1(
        sig_reg_delay1), .REG_DELAY2(sig_reg_delay2), .REG_DELAY3(
        sig_reg_delay3), .REG_DELAY4(sig_reg_delay4), .EN_IN(sig_en_dependecy), 
        .ALU_OPCODE({sig_alu_opcode[7:4], 1'b0, sig_alu_opcode[2:0]}), 
        .MUX_SEL_JAL_IMM(sig_mux_sel_jal_imm), .MUX_SEL_BIMM(sig_mux_sel_bimm), 
        .MUX_SEL_ANPC(sig_sel_anpc), .MUX_SEL_ALU_32({1'b0, 
        sig_mux_sel_alu_32[1:0]}), .MUX_SEL_ALU_1(sig_mux_sel_alu_1), 
        .ALU_OUTREG_EN(sig_alu_outreg_en), .REGBDELAY_LATCH_EN(
        sig_regbdelay_latch_en), .DRAM_WE(sig_dram_we), .LMD_LATCH_EN(
        sig_lmd_latch_en), .ALU_MA_LATCH_EN(sig_alu_ma_latch_en), .DRAM_EN(
        sig_dram_en), .MUX_SEL_WB(sig_mux_sel_wb), .RF_WE(sig_rf_we) );
  dlx_cu_FUNC_SIZE11_OP_CODE_SIZE6_CW_SIZE35 cu_0 ( .IR(sig_ir_dependency), 
        .CLK(CLK), .RST(RST), .RD1_EN(sig_rd1_en), .RD2_EN(sig_rd2_en), 
        .NPC_LATCH_DEC_EN(sig_npc_latch_dec_en), .REGA_LATCH_EN(
        sig_rega_latch_en), .REGB_LATCH_EN(sig_regb_latch_en), 
        .REGIMM_LATCH_EN(sig_regimm_latch_en), .MUX_SEL_IMM(sig_mux_sel_imm), 
        .JUMPFC(sig_jumpfc), .MUX_SEL_JAL_ADDR_LW(sig_mux_sel_jal_addr), 
        .MUX_SEL_ANPC(sig_sel_anpc), .MUX_SEL_JAL_IMM(sig_mux_sel_jal_imm), 
        .MUX_SEL_BIMM(sig_mux_sel_bimm), .ALU_OPCODE({sig_alu_opcode[7:4], 
        SYNOPSYS_UNCONNECTED__0, sig_alu_opcode[2:0]}), .MUX_SEL_ALU_32({
        SYNOPSYS_UNCONNECTED__1, sig_mux_sel_alu_32[1:0]}), .MUX_SEL_ALU_1(
        sig_mux_sel_alu_1), .ALU_OUTREG_EN(sig_alu_outreg_en), 
        .REGBDELAY_LATCH_EN(sig_regbdelay_latch_en), .DRAM_WE(sig_dram_we), 
        .LMD_LATCH_EN(sig_lmd_latch_en), .DRAM_EN(sig_dram_en), 
        .ALU_MA_LATCH_EN(sig_alu_ma_latch_en), .MUX_SEL_WB(sig_mux_sel_wb), 
        .RF_WE(sig_rf_we) );
endmodule

